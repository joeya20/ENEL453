library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

  (4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4084	)	,
(	4069	)	,
(	4055	)	,
(	4041	)	,
(	4027	)	,
(	4013	)	,
(	3999	)	,
(	3986	)	,
(	3972	)	,
(	3958	)	,
(	3945	)	,
(	3932	)	,
(	3918	)	,
(	3905	)	,
(	3892	)	,
(	3879	)	,
(	3866	)	,
(	3853	)	,
(	3840	)	,
(	3828	)	,
(	3815	)	,
(	3802	)	,
(	3790	)	,
(	3778	)	,
(	3765	)	,
(	3753	)	,
(	3741	)	,
(	3729	)	,
(	3717	)	,
(	3705	)	,
(	3693	)	,
(	3681	)	,
(	3670	)	,
(	3658	)	,
(	3646	)	,
(	3635	)	,
(	3623	)	,
(	3612	)	,
(	3601	)	,
(	3590	)	,
(	3578	)	,
(	3567	)	,
(	3556	)	,
(	3545	)	,
(	3534	)	,
(	3524	)	,
(	3513	)	,
(	3502	)	,
(	3492	)	,
(	3481	)	,
(	3470	)	,
(	3460	)	,
(	3450	)	,
(	3439	)	,
(	3429	)	,
(	3419	)	,
(	3409	)	,
(	3399	)	,
(	3389	)	,
(	3379	)	,
(	3369	)	,
(	3359	)	,
(	3349	)	,
(	3339	)	,
(	3330	)	,
(	3320	)	,
(	3310	)	,
(	3301	)	,
(	3291	)	,
(	3282	)	,
(	3272	)	,
(	3263	)	,
(	3254	)	,
(	3245	)	,
(	3235	)	,
(	3226	)	,
(	3217	)	,
(	3208	)	,
(	3199	)	,
(	3190	)	,
(	3181	)	,
(	3173	)	,
(	3164	)	,
(	3155	)	,
(	3146	)	,
(	3138	)	,
(	3129	)	,
(	3121	)	,
(	3112	)	,
(	3104	)	,
(	3095	)	,
(	3087	)	,
(	3078	)	,
(	3070	)	,
(	3062	)	,
(	3054	)	,
(	3045	)	,
(	3037	)	,
(	3029	)	,
(	3021	)	,
(	3013	)	,
(	3005	)	,
(	2997	)	,
(	2989	)	,
(	2982	)	,
(	2974	)	,
(	2966	)	,
(	2958	)	,
(	2951	)	,
(	2943	)	,
(	2935	)	,
(	2928	)	,
(	2920	)	,
(	2913	)	,
(	2905	)	,
(	2898	)	,
(	2891	)	,
(	2883	)	,
(	2876	)	,
(	2869	)	,
(	2861	)	,
(	2854	)	,
(	2847	)	,
(	2840	)	,
(	2833	)	,
(	2826	)	,
(	2819	)	,
(	2812	)	,
(	2805	)	,
(	2798	)	,
(	2791	)	,
(	2784	)	,
(	2777	)	,
(	2770	)	,
(	2764	)	,
(	2757	)	,
(	2750	)	,
(	2744	)	,
(	2737	)	,
(	2730	)	,
(	2724	)	,
(	2717	)	,
(	2711	)	,
(	2704	)	,
(	2698	)	,
(	2691	)	,
(	2685	)	,
(	2679	)	,
(	2672	)	,
(	2666	)	,
(	2660	)	,
(	2653	)	,
(	2647	)	,
(	2641	)	,
(	2635	)	,
(	2629	)	,
(	2622	)	,
(	2616	)	,
(	2610	)	,
(	2604	)	,
(	2598	)	,
(	2592	)	,
(	2586	)	,
(	2580	)	,
(	2575	)	,
(	2569	)	,
(	2563	)	,
(	2557	)	,
(	2551	)	,
(	2545	)	,
(	2540	)	,
(	2534	)	,
(	2528	)	,
(	2523	)	,
(	2517	)	,
(	2511	)	,
(	2506	)	,
(	2500	)	,
(	2495	)	,
(	2489	)	,
(	2484	)	,
(	2478	)	,
(	2473	)	,
(	2467	)	,
(	2462	)	,
(	2456	)	,
(	2451	)	,
(	2446	)	,
(	2440	)	,
(	2435	)	,
(	2430	)	,
(	2424	)	,
(	2419	)	,
(	2414	)	,
(	2409	)	,
(	2404	)	,
(	2399	)	,
(	2393	)	,
(	2388	)	,
(	2383	)	,
(	2378	)	,
(	2373	)	,
(	2368	)	,
(	2363	)	,
(	2358	)	,
(	2353	)	,
(	2348	)	,
(	2343	)	,
(	2338	)	,
(	2333	)	,
(	2329	)	,
(	2324	)	,
(	2319	)	,
(	2314	)	,
(	2309	)	,
(	2305	)	,
(	2300	)	,
(	2295	)	,
(	2290	)	,
(	2286	)	,
(	2281	)	,
(	2276	)	,
(	2272	)	,
(	2267	)	,
(	2263	)	,
(	2258	)	,
(	2253	)	,
(	2249	)	,
(	2244	)	,
(	2240	)	,
(	2235	)	,
(	2231	)	,
(	2226	)	,
(	2222	)	,
(	2218	)	,
(	2213	)	,
(	2209	)	,
(	2204	)	,
(	2200	)	,
(	2196	)	,
(	2191	)	,
(	2187	)	,
(	2183	)	,
(	2179	)	,
(	2174	)	,
(	2170	)	,
(	2166	)	,
(	2162	)	,
(	2157	)	,
(	2153	)	,
(	2149	)	,
(	2145	)	,
(	2141	)	,
(	2137	)	,
(	2133	)	,
(	2128	)	,
(	2124	)	,
(	2120	)	,
(	2116	)	,
(	2112	)	,
(	2108	)	,
(	2104	)	,
(	2100	)	,
(	2096	)	,
(	2092	)	,
(	2088	)	,
(	2084	)	,
(	2081	)	,
(	2077	)	,
(	2073	)	,
(	2069	)	,
(	2065	)	,
(	2061	)	,
(	2057	)	,
(	2054	)	,
(	2050	)	,
(	2046	)	,
(	2042	)	,
(	2038	)	,
(	2035	)	,
(	2031	)	,
(	2027	)	,
(	2024	)	,
(	2020	)	,
(	2016	)	,
(	2013	)	,
(	2009	)	,
(	2005	)	,
(	2002	)	,
(	1998	)	,
(	1994	)	,
(	1991	)	,
(	1987	)	,
(	1984	)	,
(	1980	)	,
(	1977	)	,
(	1973	)	,
(	1970	)	,
(	1966	)	,
(	1963	)	,
(	1959	)	,
(	1956	)	,
(	1952	)	,
(	1949	)	,
(	1945	)	,
(	1942	)	,
(	1938	)	,
(	1935	)	,
(	1932	)	,
(	1928	)	,
(	1925	)	,
(	1922	)	,
(	1918	)	,
(	1915	)	,
(	1912	)	,
(	1908	)	,
(	1905	)	,
(	1902	)	,
(	1898	)	,
(	1895	)	,
(	1892	)	,
(	1889	)	,
(	1885	)	,
(	1882	)	,
(	1879	)	,
(	1876	)	,
(	1873	)	,
(	1869	)	,
(	1866	)	,
(	1863	)	,
(	1860	)	,
(	1857	)	,
(	1854	)	,
(	1850	)	,
(	1847	)	,
(	1844	)	,
(	1841	)	,
(	1838	)	,
(	1835	)	,
(	1832	)	,
(	1829	)	,
(	1826	)	,
(	1823	)	,
(	1820	)	,
(	1817	)	,
(	1814	)	,
(	1811	)	,
(	1808	)	,
(	1805	)	,
(	1802	)	,
(	1799	)	,
(	1796	)	,
(	1793	)	,
(	1790	)	,
(	1787	)	,
(	1784	)	,
(	1781	)	,
(	1779	)	,
(	1776	)	,
(	1773	)	,
(	1770	)	,
(	1767	)	,
(	1764	)	,
(	1761	)	,
(	1759	)	,
(	1756	)	,
(	1753	)	,
(	1750	)	,
(	1747	)	,
(	1745	)	,
(	1742	)	,
(	1739	)	,
(	1736	)	,
(	1734	)	,
(	1731	)	,
(	1728	)	,
(	1725	)	,
(	1723	)	,
(	1720	)	,
(	1717	)	,
(	1715	)	,
(	1712	)	,
(	1709	)	,
(	1707	)	,
(	1704	)	,
(	1701	)	,
(	1699	)	,
(	1696	)	,
(	1693	)	,
(	1691	)	,
(	1688	)	,
(	1685	)	,
(	1683	)	,
(	1680	)	,
(	1678	)	,
(	1675	)	,
(	1673	)	,
(	1670	)	,
(	1667	)	,
(	1665	)	,
(	1662	)	,
(	1660	)	,
(	1657	)	,
(	1655	)	,
(	1652	)	,
(	1650	)	,
(	1647	)	,
(	1645	)	,
(	1642	)	,
(	1640	)	,
(	1637	)	,
(	1635	)	,
(	1633	)	,
(	1630	)	,
(	1628	)	,
(	1625	)	,
(	1623	)	,
(	1620	)	,
(	1618	)	,
(	1616	)	,
(	1613	)	,
(	1611	)	,
(	1608	)	,
(	1606	)	,
(	1604	)	,
(	1601	)	,
(	1599	)	,
(	1597	)	,
(	1594	)	,
(	1592	)	,
(	1590	)	,
(	1587	)	,
(	1585	)	,
(	1583	)	,
(	1580	)	,
(	1578	)	,
(	1576	)	,
(	1574	)	,
(	1571	)	,
(	1569	)	,
(	1567	)	,
(	1565	)	,
(	1562	)	,
(	1560	)	,
(	1558	)	,
(	1556	)	,
(	1553	)	,
(	1551	)	,
(	1549	)	,
(	1547	)	,
(	1544	)	,
(	1542	)	,
(	1540	)	,
(	1538	)	,
(	1536	)	,
(	1534	)	,
(	1531	)	,
(	1529	)	,
(	1527	)	,
(	1525	)	,
(	1523	)	,
(	1521	)	,
(	1519	)	,
(	1516	)	,
(	1514	)	,
(	1512	)	,
(	1510	)	,
(	1508	)	,
(	1506	)	,
(	1504	)	,
(	1502	)	,
(	1500	)	,
(	1498	)	,
(	1496	)	,
(	1493	)	,
(	1491	)	,
(	1489	)	,
(	1487	)	,
(	1485	)	,
(	1483	)	,
(	1481	)	,
(	1479	)	,
(	1477	)	,
(	1475	)	,
(	1473	)	,
(	1471	)	,
(	1469	)	,
(	1467	)	,
(	1465	)	,
(	1463	)	,
(	1461	)	,
(	1459	)	,
(	1457	)	,
(	1455	)	,
(	1453	)	,
(	1451	)	,
(	1449	)	,
(	1448	)	,
(	1446	)	,
(	1444	)	,
(	1442	)	,
(	1440	)	,
(	1438	)	,
(	1436	)	,
(	1434	)	,
(	1432	)	,
(	1430	)	,
(	1428	)	,
(	1427	)	,
(	1425	)	,
(	1423	)	,
(	1421	)	,
(	1419	)	,
(	1417	)	,
(	1415	)	,
(	1413	)	,
(	1412	)	,
(	1410	)	,
(	1408	)	,
(	1406	)	,
(	1404	)	,
(	1402	)	,
(	1401	)	,
(	1399	)	,
(	1397	)	,
(	1395	)	,
(	1393	)	,
(	1392	)	,
(	1390	)	,
(	1388	)	,
(	1386	)	,
(	1384	)	,
(	1383	)	,
(	1381	)	,
(	1379	)	,
(	1377	)	,
(	1376	)	,
(	1374	)	,
(	1372	)	,
(	1370	)	,
(	1369	)	,
(	1367	)	,
(	1365	)	,
(	1363	)	,
(	1362	)	,
(	1360	)	,
(	1358	)	,
(	1357	)	,
(	1355	)	,
(	1353	)	,
(	1351	)	,
(	1350	)	,
(	1348	)	,
(	1346	)	,
(	1345	)	,
(	1343	)	,
(	1341	)	,
(	1340	)	,
(	1338	)	,
(	1336	)	,
(	1335	)	,
(	1333	)	,
(	1331	)	,
(	1330	)	,
(	1328	)	,
(	1326	)	,
(	1325	)	,
(	1323	)	,
(	1322	)	,
(	1320	)	,
(	1318	)	,
(	1317	)	,
(	1315	)	,
(	1313	)	,
(	1312	)	,
(	1310	)	,
(	1309	)	,
(	1307	)	,
(	1305	)	,
(	1304	)	,
(	1302	)	,
(	1301	)	,
(	1299	)	,
(	1298	)	,
(	1296	)	,
(	1294	)	,
(	1293	)	,
(	1291	)	,
(	1290	)	,
(	1288	)	,
(	1287	)	,
(	1285	)	,
(	1284	)	,
(	1282	)	,
(	1281	)	,
(	1279	)	,
(	1277	)	,
(	1276	)	,
(	1274	)	,
(	1273	)	,
(	1271	)	,
(	1270	)	,
(	1268	)	,
(	1267	)	,
(	1265	)	,
(	1264	)	,
(	1262	)	,
(	1261	)	,
(	1259	)	,
(	1258	)	,
(	1256	)	,
(	1255	)	,
(	1254	)	,
(	1252	)	,
(	1251	)	,
(	1249	)	,
(	1248	)	,
(	1246	)	,
(	1245	)	,
(	1243	)	,
(	1242	)	,
(	1240	)	,
(	1239	)	,
(	1238	)	,
(	1236	)	,
(	1235	)	,
(	1233	)	,
(	1232	)	,
(	1230	)	,
(	1229	)	,
(	1228	)	,
(	1226	)	,
(	1225	)	,
(	1223	)	,
(	1222	)	,
(	1221	)	,
(	1219	)	,
(	1218	)	,
(	1216	)	,
(	1215	)	,
(	1214	)	,
(	1212	)	,
(	1211	)	,
(	1210	)	,
(	1208	)	,
(	1207	)	,
(	1205	)	,
(	1204	)	,
(	1203	)	,
(	1201	)	,
(	1200	)	,
(	1199	)	,
(	1197	)	,
(	1196	)	,
(	1195	)	,
(	1193	)	,
(	1192	)	,
(	1191	)	,
(	1189	)	,
(	1188	)	,
(	1187	)	,
(	1185	)	,
(	1184	)	,
(	1183	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1178	)	,
(	1176	)	,
(	1175	)	,
(	1174	)	,
(	1172	)	,
(	1171	)	,
(	1170	)	,
(	1169	)	,
(	1167	)	,
(	1166	)	,
(	1165	)	,
(	1163	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1158	)	,
(	1157	)	,
(	1156	)	,
(	1155	)	,
(	1153	)	,
(	1152	)	,
(	1151	)	,
(	1150	)	,
(	1148	)	,
(	1147	)	,
(	1146	)	,
(	1145	)	,
(	1143	)	,
(	1142	)	,
(	1141	)	,
(	1140	)	,
(	1139	)	,
(	1137	)	,
(	1136	)	,
(	1135	)	,
(	1134	)	,
(	1132	)	,
(	1131	)	,
(	1130	)	,
(	1129	)	,
(	1128	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1116	)	,
(	1115	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1108	)	,
(	1106	)	,
(	1105	)	,
(	1104	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1098	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1067	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1052	)	,
(	1051	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1025	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1005	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	989	)	,
(	989	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	977	)	,
(	977	)	,
(	976	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	972	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	968	)	,
(	968	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	962	)	,
(	961	)	,
(	961	)	,
(	960	)	,
(	959	)	,
(	958	)	,
(	957	)	,
(	956	)	,
(	955	)	,
(	954	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	951	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	948	)	,
(	947	)	,
(	946	)	,
(	945	)	,
(	944	)	,
(	943	)	,
(	942	)	,
(	942	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	938	)	,
(	937	)	,
(	937	)	,
(	936	)	,
(	935	)	,
(	934	)	,
(	933	)	,
(	932	)	,
(	932	)	,
(	931	)	,
(	930	)	,
(	929	)	,
(	928	)	,
(	927	)	,
(	927	)	,
(	926	)	,
(	925	)	,
(	924	)	,
(	923	)	,
(	923	)	,
(	922	)	,
(	921	)	,
(	920	)	,
(	919	)	,
(	918	)	,
(	918	)	,
(	917	)	,
(	916	)	,
(	915	)	,
(	914	)	,
(	914	)	,
(	913	)	,
(	912	)	,
(	911	)	,
(	910	)	,
(	910	)	,
(	909	)	,
(	908	)	,
(	907	)	,
(	907	)	,
(	906	)	,
(	905	)	,
(	904	)	,
(	903	)	,
(	903	)	,
(	902	)	,
(	901	)	,
(	900	)	,
(	900	)	,
(	899	)	,
(	898	)	,
(	897	)	,
(	896	)	,
(	896	)	,
(	895	)	,
(	894	)	,
(	893	)	,
(	893	)	,
(	892	)	,
(	891	)	,
(	890	)	,
(	890	)	,
(	889	)	,
(	888	)	,
(	887	)	,
(	887	)	,
(	886	)	,
(	885	)	,
(	884	)	,
(	884	)	,
(	883	)	,
(	882	)	,
(	881	)	,
(	881	)	,
(	880	)	,
(	879	)	,
(	878	)	,
(	878	)	,
(	877	)	,
(	876	)	,
(	875	)	,
(	875	)	,
(	874	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	868	)	,
(	867	)	,
(	867	)	,
(	866	)	,
(	865	)	,
(	865	)	,
(	864	)	,
(	863	)	,
(	862	)	,
(	862	)	,
(	861	)	,
(	860	)	,
(	860	)	,
(	859	)	,
(	858	)	,
(	857	)	,
(	857	)	,
(	856	)	,
(	855	)	,
(	855	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	851	)	,
(	850	)	,
(	850	)	,
(	849	)	,
(	848	)	,
(	848	)	,
(	847	)	,
(	846	)	,
(	846	)	,
(	845	)	,
(	844	)	,
(	844	)	,
(	843	)	,
(	842	)	,
(	842	)	,
(	841	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	837	)	,
(	837	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	833	)	,
(	833	)	,
(	832	)	,
(	831	)	,
(	831	)	,
(	830	)	,
(	829	)	,
(	829	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	824	)	,
(	823	)	,
(	822	)	,
(	822	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	816	)	,
(	816	)	,
(	815	)	,
(	814	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	811	)	,
(	811	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	808	)	,
(	807	)	,
(	806	)	,
(	806	)	,
(	805	)	,
(	804	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	796	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	793	)	,
(	793	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	769	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	755	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	747	)	,
(	747	)	,
(	746	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	742	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	729	)	,
(	729	)	,
(	728	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	700	)	,
(	699	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	697	)	,
(	696	)	,
(	696	)	,
(	695	)	,
(	695	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	684	)	,
(	683	)	,
(	683	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	674	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	667	)	,
(	667	)	,
(	666	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	664	)	,
(	664	)	,
(	663	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	661	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	658	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	655	)	,
(	655	)	,
(	654	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	650	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	647	)	,
(	646	)	,
(	646	)	,
(	646	)	,
(	645	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	643	)	,
(	643	)	,
(	642	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	639	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	637	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	635	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	622	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	619	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	617	)	,
(	617	)	,
(	616	)	,
(	616	)	,
(	616	)	,
(	615	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	613	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	610	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	608	)	,
(	607	)	,
(	607	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	601	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	596	)	,
(	596	)	,
(	595	)	,
(	595	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	592	)	,
(	592	)	,
(	591	)	,
(	591	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	586	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	584	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	582	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	579	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	577	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	574	)	,
(	574	)	,
(	574	)	,
(	573	)	,
(	573	)	,
(	573	)	,
(	572	)	,
(	572	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	570	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	567	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	564	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	561	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	559	)	,
(	559	)	,
(	558	)	,
(	558	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	551	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	548	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	539	)	,
(	539	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	537	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	

);

--Eqn 50,000,000/ (4096*(49/4)-(9x/1600))
--Where x is the distance ranging from 400 mm to 2000mm
-- x<=400mm then the period = 50,000,000/(4096 * 10Hz))  
-- x>=2000mm then the period = 50,000,000/(4096 * 1Hz))  
constant d27seg_LUT : array_1d := (
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 610 ),
( 626 ),
( 627 ),
( 627 ),
( 627 ),
( 628 ),
( 628 ),
( 629 ),
( 629 ),
( 629 ),
( 630 ),
( 630 ),
( 630 ),
( 631 ),
( 631 ),
( 631 ),
( 632 ),
( 632 ),
( 633 ),
( 633 ),
( 633 ),
( 634 ),
( 634 ),
( 634 ),
( 635 ),
( 635 ),
( 636 ),
( 636 ),
( 636 ),
( 637 ),
( 637 ),
( 637 ),
( 638 ),
( 638 ),
( 639 ),
( 639 ),
( 639 ),
( 640 ),
( 640 ),
( 640 ),
( 641 ),
( 641 ),
( 642 ),
( 642 ),
( 642 ),
( 643 ),
( 643 ),
( 643 ),
( 644 ),
( 644 ),
( 645 ),
( 645 ),
( 645 ),
( 646 ),
( 646 ),
( 647 ),
( 647 ),
( 647 ),
( 648 ),
( 648 ),
( 648 ),
( 649 ),
( 649 ),
( 650 ),
( 650 ),
( 650 ),
( 651 ),
( 651 ),
( 652 ),
( 652 ),
( 652 ),
( 653 ),
( 653 ),
( 654 ),
( 654 ),
( 654 ),
( 655 ),
( 655 ),
( 655 ),
( 656 ),
( 656 ),
( 657 ),
( 657 ),
( 657 ),
( 658 ),
( 658 ),
( 659 ),
( 659 ),
( 659 ),
( 660 ),
( 660 ),
( 661 ),
( 661 ),
( 661 ),
( 662 ),
( 662 ),
( 663 ),
( 663 ),
( 664 ),
( 664 ),
( 664 ),
( 665 ),
( 665 ),
( 666 ),
( 666 ),
( 666 ),
( 667 ),
( 667 ),
( 668 ),
( 668 ),
( 668 ),
( 669 ),
( 669 ),
( 670 ),
( 670 ),
( 670 ),
( 671 ),
( 671 ),
( 672 ),
( 672 ),
( 673 ),
( 673 ),
( 673 ),
( 674 ),
( 674 ),
( 675 ),
( 675 ),
( 675 ),
( 676 ),
( 676 ),
( 677 ),
( 677 ),
( 678 ),
( 678 ),
( 678 ),
( 679 ),
( 679 ),
( 680 ),
( 680 ),
( 681 ),
( 681 ),
( 681 ),
( 682 ),
( 682 ),
( 683 ),
( 683 ),
( 684 ),
( 684 ),
( 684 ),
( 685 ),
( 685 ),
( 686 ),
( 686 ),
( 687 ),
( 687 ),
( 687 ),
( 688 ),
( 688 ),
( 689 ),
( 689 ),
( 690 ),
( 690 ),
( 691 ),
( 691 ),
( 691 ),
( 692 ),
( 692 ),
( 693 ),
( 693 ),
( 694 ),
( 694 ),
( 695 ),
( 695 ),
( 695 ),
( 696 ),
( 696 ),
( 697 ),
( 697 ),
( 698 ),
( 698 ),
( 699 ),
( 699 ),
( 699 ),
( 700 ),
( 700 ),
( 701 ),
( 701 ),
( 702 ),
( 702 ),
( 703 ),
( 703 ),
( 704 ),
( 704 ),
( 704 ),
( 705 ),
( 705 ),
( 706 ),
( 706 ),
( 707 ),
( 707 ),
( 708 ),
( 708 ),
( 709 ),
( 709 ),
( 710 ),
( 710 ),
( 710 ),
( 711 ),
( 711 ),
( 712 ),
( 712 ),
( 713 ),
( 713 ),
( 714 ),
( 714 ),
( 715 ),
( 715 ),
( 716 ),
( 716 ),
( 717 ),
( 717 ),
( 717 ),
( 718 ),
( 718 ),
( 719 ),
( 719 ),
( 720 ),
( 720 ),
( 721 ),
( 721 ),
( 722 ),
( 722 ),
( 723 ),
( 723 ),
( 724 ),
( 724 ),
( 725 ),
( 725 ),
( 726 ),
( 726 ),
( 727 ),
( 727 ),
( 728 ),
( 728 ),
( 729 ),
( 729 ),
( 730 ),
( 730 ),
( 731 ),
( 731 ),
( 732 ),
( 732 ),
( 732 ),
( 733 ),
( 733 ),
( 734 ),
( 734 ),
( 735 ),
( 735 ),
( 736 ),
( 736 ),
( 737 ),
( 737 ),
( 738 ),
( 738 ),
( 739 ),
( 739 ),
( 740 ),
( 740 ),
( 741 ),
( 742 ),
( 742 ),
( 743 ),
( 743 ),
( 744 ),
( 744 ),
( 745 ),
( 745 ),
( 746 ),
( 746 ),
( 747 ),
( 747 ),
( 748 ),
( 748 ),
( 749 ),
( 749 ),
( 750 ),
( 750 ),
( 751 ),
( 751 ),
( 752 ),
( 752 ),
( 753 ),
( 753 ),
( 754 ),
( 754 ),
( 755 ),
( 755 ),
( 756 ),
( 756 ),
( 757 ),
( 758 ),
( 758 ),
( 759 ),
( 759 ),
( 760 ),
( 760 ),
( 761 ),
( 761 ),
( 762 ),
( 762 ),
( 763 ),
( 763 ),
( 764 ),
( 764 ),
( 765 ),
( 766 ),
( 766 ),
( 767 ),
( 767 ),
( 768 ),
( 768 ),
( 769 ),
( 769 ),
( 770 ),
( 770 ),
( 771 ),
( 772 ),
( 772 ),
( 773 ),
( 773 ),
( 774 ),
( 774 ),
( 775 ),
( 775 ),
( 776 ),
( 777 ),
( 777 ),
( 778 ),
( 778 ),
( 779 ),
( 779 ),
( 780 ),
( 780 ),
( 781 ),
( 782 ),
( 782 ),
( 783 ),
( 783 ),
( 784 ),
( 784 ),
( 785 ),
( 786 ),
( 786 ),
( 787 ),
( 787 ),
( 788 ),
( 788 ),
( 789 ),
( 790 ),
( 790 ),
( 791 ),
( 791 ),
( 792 ),
( 792 ),
( 793 ),
( 794 ),
( 794 ),
( 795 ),
( 795 ),
( 796 ),
( 796 ),
( 797 ),
( 798 ),
( 798 ),
( 799 ),
( 799 ),
( 800 ),
( 801 ),
( 801 ),
( 802 ),
( 802 ),
( 803 ),
( 804 ),
( 804 ),
( 805 ),
( 805 ),
( 806 ),
( 807 ),
( 807 ),
( 808 ),
( 808 ),
( 809 ),
( 810 ),
( 810 ),
( 811 ),
( 811 ),
( 812 ),
( 813 ),
( 813 ),
( 814 ),
( 814 ),
( 815 ),
( 816 ),
( 816 ),
( 817 ),
( 817 ),
( 818 ),
( 819 ),
( 819 ),
( 820 ),
( 821 ),
( 821 ),
( 822 ),
( 822 ),
( 823 ),
( 824 ),
( 824 ),
( 825 ),
( 826 ),
( 826 ),
( 827 ),
( 827 ),
( 828 ),
( 829 ),
( 829 ),
( 830 ),
( 831 ),
( 831 ),
( 832 ),
( 833 ),
( 833 ),
( 834 ),
( 834 ),
( 835 ),
( 836 ),
( 836 ),
( 837 ),
( 838 ),
( 838 ),
( 839 ),
( 840 ),
( 840 ),
( 841 ),
( 842 ),
( 842 ),
( 843 ),
( 844 ),
( 844 ),
( 845 ),
( 846 ),
( 846 ),
( 847 ),
( 847 ),
( 848 ),
( 849 ),
( 849 ),
( 850 ),
( 851 ),
( 851 ),
( 852 ),
( 853 ),
( 853 ),
( 854 ),
( 855 ),
( 856 ),
( 856 ),
( 857 ),
( 858 ),
( 858 ),
( 859 ),
( 860 ),
( 860 ),
( 861 ),
( 862 ),
( 862 ),
( 863 ),
( 864 ),
( 864 ),
( 865 ),
( 866 ),
( 866 ),
( 867 ),
( 868 ),
( 869 ),
( 869 ),
( 870 ),
( 871 ),
( 871 ),
( 872 ),
( 873 ),
( 873 ),
( 874 ),
( 875 ),
( 876 ),
( 876 ),
( 877 ),
( 878 ),
( 878 ),
( 879 ),
( 880 ),
( 880 ),
( 881 ),
( 882 ),
( 883 ),
( 883 ),
( 884 ),
( 885 ),
( 886 ),
( 886 ),
( 887 ),
( 888 ),
( 888 ),
( 889 ),
( 890 ),
( 891 ),
( 891 ),
( 892 ),
( 893 ),
( 894 ),
( 894 ),
( 895 ),
( 896 ),
( 897 ),
( 897 ),
( 898 ),
( 899 ),
( 899 ),
( 900 ),
( 901 ),
( 902 ),
( 902 ),
( 903 ),
( 904 ),
( 905 ),
( 905 ),
( 906 ),
( 907 ),
( 908 ),
( 909 ),
( 909 ),
( 910 ),
( 911 ),
( 912 ),
( 912 ),
( 913 ),
( 914 ),
( 915 ),
( 915 ),
( 916 ),
( 917 ),
( 918 ),
( 919 ),
( 919 ),
( 920 ),
( 921 ),
( 922 ),
( 922 ),
( 923 ),
( 924 ),
( 925 ),
( 926 ),
( 926 ),
( 927 ),
( 928 ),
( 929 ),
( 930 ),
( 930 ),
( 931 ),
( 932 ),
( 933 ),
( 934 ),
( 934 ),
( 935 ),
( 936 ),
( 937 ),
( 938 ),
( 938 ),
( 939 ),
( 940 ),
( 941 ),
( 942 ),
( 942 ),
( 943 ),
( 944 ),
( 945 ),
( 946 ),
( 947 ),
( 947 ),
( 948 ),
( 949 ),
( 950 ),
( 951 ),
( 952 ),
( 952 ),
( 953 ),
( 954 ),
( 955 ),
( 956 ),
( 957 ),
( 957 ),
( 958 ),
( 959 ),
( 960 ),
( 961 ),
( 962 ),
( 963 ),
( 963 ),
( 964 ),
( 965 ),
( 966 ),
( 967 ),
( 968 ),
( 969 ),
( 969 ),
( 970 ),
( 971 ),
( 972 ),
( 973 ),
( 974 ),
( 975 ),
( 975 ),
( 976 ),
( 977 ),
( 978 ),
( 979 ),
( 980 ),
( 981 ),
( 982 ),
( 983 ),
( 983 ),
( 984 ),
( 985 ),
( 986 ),
( 987 ),
( 988 ),
( 989 ),
( 990 ),
( 991 ),
( 992 ),
( 992 ),
( 993 ),
( 994 ),
( 995 ),
( 996 ),
( 997 ),
( 998 ),
( 999 ),
( 1000 ),
( 1001 ),
( 1002 ),
( 1003 ),
( 1003 ),
( 1004 ),
( 1005 ),
( 1006 ),
( 1007 ),
( 1008 ),
( 1009 ),
( 1010 ),
( 1011 ),
( 1012 ),
( 1013 ),
( 1014 ),
( 1015 ),
( 1016 ),
( 1017 ),
( 1018 ),
( 1019 ),
( 1019 ),
( 1020 ),
( 1021 ),
( 1022 ),
( 1023 ),
( 1024 ),
( 1025 ),
( 1026 ),
( 1027 ),
( 1028 ),
( 1029 ),
( 1030 ),
( 1031 ),
( 1032 ),
( 1033 ),
( 1034 ),
( 1035 ),
( 1036 ),
( 1037 ),
( 1038 ),
( 1039 ),
( 1040 ),
( 1041 ),
( 1042 ),
( 1043 ),
( 1044 ),
( 1045 ),
( 1046 ),
( 1047 ),
( 1048 ),
( 1049 ),
( 1050 ),
( 1051 ),
( 1052 ),
( 1053 ),
( 1054 ),
( 1055 ),
( 1056 ),
( 1057 ),
( 1058 ),
( 1059 ),
( 1060 ),
( 1061 ),
( 1062 ),
( 1063 ),
( 1064 ),
( 1066 ),
( 1067 ),
( 1068 ),
( 1069 ),
( 1070 ),
( 1071 ),
( 1072 ),
( 1073 ),
( 1074 ),
( 1075 ),
( 1076 ),
( 1077 ),
( 1078 ),
( 1079 ),
( 1080 ),
( 1081 ),
( 1083 ),
( 1084 ),
( 1085 ),
( 1086 ),
( 1087 ),
( 1088 ),
( 1089 ),
( 1090 ),
( 1091 ),
( 1092 ),
( 1093 ),
( 1095 ),
( 1096 ),
( 1097 ),
( 1098 ),
( 1099 ),
( 1100 ),
( 1101 ),
( 1102 ),
( 1103 ),
( 1105 ),
( 1106 ),
( 1107 ),
( 1108 ),
( 1109 ),
( 1110 ),
( 1111 ),
( 1113 ),
( 1114 ),
( 1115 ),
( 1116 ),
( 1117 ),
( 1118 ),
( 1119 ),
( 1121 ),
( 1122 ),
( 1123 ),
( 1124 ),
( 1125 ),
( 1126 ),
( 1128 ),
( 1129 ),
( 1130 ),
( 1131 ),
( 1132 ),
( 1133 ),
( 1135 ),
( 1136 ),
( 1137 ),
( 1138 ),
( 1139 ),
( 1141 ),
( 1142 ),
( 1143 ),
( 1144 ),
( 1145 ),
( 1147 ),
( 1148 ),
( 1149 ),
( 1150 ),
( 1151 ),
( 1153 ),
( 1154 ),
( 1155 ),
( 1156 ),
( 1158 ),
( 1159 ),
( 1160 ),
( 1161 ),
( 1163 ),
( 1164 ),
( 1165 ),
( 1166 ),
( 1168 ),
( 1169 ),
( 1170 ),
( 1171 ),
( 1173 ),
( 1174 ),
( 1175 ),
( 1176 ),
( 1178 ),
( 1179 ),
( 1180 ),
( 1182 ),
( 1183 ),
( 1184 ),
( 1185 ),
( 1187 ),
( 1188 ),
( 1189 ),
( 1191 ),
( 1192 ),
( 1193 ),
( 1195 ),
( 1196 ),
( 1197 ),
( 1199 ),
( 1200 ),
( 1201 ),
( 1203 ),
( 1204 ),
( 1205 ),
( 1207 ),
( 1208 ),
( 1209 ),
( 1211 ),
( 1212 ),
( 1213 ),
( 1215 ),
( 1216 ),
( 1217 ),
( 1219 ),
( 1220 ),
( 1221 ),
( 1223 ),
( 1224 ),
( 1226 ),
( 1227 ),
( 1228 ),
( 1230 ),
( 1231 ),
( 1233 ),
( 1234 ),
( 1235 ),
( 1237 ),
( 1238 ),
( 1240 ),
( 1241 ),
( 1242 ),
( 1244 ),
( 1245 ),
( 1247 ),
( 1248 ),
( 1250 ),
( 1251 ),
( 1252 ),
( 1254 ),
( 1255 ),
( 1257 ),
( 1258 ),
( 1260 ),
( 1261 ),
( 1263 ),
( 1264 ),
( 1266 ),
( 1267 ),
( 1269 ),
( 1270 ),
( 1272 ),
( 1273 ),
( 1275 ),
( 1276 ),
( 1278 ),
( 1279 ),
( 1281 ),
( 1282 ),
( 1284 ),
( 1285 ),
( 1287 ),
( 1288 ),
( 1290 ),
( 1291 ),
( 1293 ),
( 1294 ),
( 1296 ),
( 1297 ),
( 1299 ),
( 1301 ),
( 1302 ),
( 1304 ),
( 1305 ),
( 1307 ),
( 1308 ),
( 1310 ),
( 1312 ),
( 1313 ),
( 1315 ),
( 1316 ),
( 1318 ),
( 1320 ),
( 1321 ),
( 1323 ),
( 1324 ),
( 1326 ),
( 1328 ),
( 1329 ),
( 1331 ),
( 1332 ),
( 1334 ),
( 1336 ),
( 1337 ),
( 1339 ),
( 1341 ),
( 1342 ),
( 1344 ),
( 1346 ),
( 1347 ),
( 1349 ),
( 1351 ),
( 1352 ),
( 1354 ),
( 1356 ),
( 1357 ),
( 1359 ),
( 1361 ),
( 1363 ),
( 1364 ),
( 1366 ),
( 1368 ),
( 1369 ),
( 1371 ),
( 1373 ),
( 1375 ),
( 1376 ),
( 1378 ),
( 1380 ),
( 1382 ),
( 1383 ),
( 1385 ),
( 1387 ),
( 1389 ),
( 1391 ),
( 1392 ),
( 1394 ),
( 1396 ),
( 1398 ),
( 1399 ),
( 1401 ),
( 1403 ),
( 1405 ),
( 1407 ),
( 1409 ),
( 1410 ),
( 1412 ),
( 1414 ),
( 1416 ),
( 1418 ),
( 1420 ),
( 1421 ),
( 1423 ),
( 1425 ),
( 1427 ),
( 1429 ),
( 1431 ),
( 1433 ),
( 1435 ),
( 1437 ),
( 1438 ),
( 1440 ),
( 1442 ),
( 1444 ),
( 1446 ),
( 1448 ),
( 1450 ),
( 1452 ),
( 1454 ),
( 1456 ),
( 1458 ),
( 1460 ),
( 1462 ),
( 1464 ),
( 1466 ),
( 1468 ),
( 1470 ),
( 1472 ),
( 1474 ),
( 1476 ),
( 1478 ),
( 1480 ),
( 1482 ),
( 1484 ),
( 1486 ),
( 1488 ),
( 1490 ),
( 1492 ),
( 1494 ),
( 1496 ),
( 1498 ),
( 1500 ),
( 1502 ),
( 1504 ),
( 1506 ),
( 1508 ),
( 1511 ),
( 1513 ),
( 1515 ),
( 1517 ),
( 1519 ),
( 1521 ),
( 1523 ),
( 1525 ),
( 1528 ),
( 1530 ),
( 1532 ),
( 1534 ),
( 1536 ),
( 1538 ),
( 1541 ),
( 1543 ),
( 1545 ),
( 1547 ),
( 1549 ),
( 1552 ),
( 1554 ),
( 1556 ),
( 1558 ),
( 1561 ),
( 1563 ),
( 1565 ),
( 1567 ),
( 1570 ),
( 1572 ),
( 1574 ),
( 1576 ),
( 1579 ),
( 1581 ),
( 1583 ),
( 1586 ),
( 1588 ),
( 1590 ),
( 1593 ),
( 1595 ),
( 1597 ),
( 1600 ),
( 1602 ),
( 1604 ),
( 1607 ),
( 1609 ),
( 1611 ),
( 1614 ),
( 1616 ),
( 1619 ),
( 1621 ),
( 1624 ),
( 1626 ),
( 1628 ),
( 1631 ),
( 1633 ),
( 1636 ),
( 1638 ),
( 1641 ),
( 1643 ),
( 1646 ),
( 1648 ),
( 1651 ),
( 1653 ),
( 1656 ),
( 1658 ),
( 1661 ),
( 1663 ),
( 1666 ),
( 1668 ),
( 1671 ),
( 1674 ),
( 1676 ),
( 1679 ),
( 1681 ),
( 1684 ),
( 1687 ),
( 1689 ),
( 1692 ),
( 1695 ),
( 1697 ),
( 1700 ),
( 1703 ),
( 1705 ),
( 1708 ),
( 1711 ),
( 1713 ),
( 1716 ),
( 1719 ),
( 1721 ),
( 1724 ),
( 1727 ),
( 1730 ),
( 1732 ),
( 1735 ),
( 1738 ),
( 1741 ),
( 1744 ),
( 1746 ),
( 1749 ),
( 1752 ),
( 1755 ),
( 1758 ),
( 1761 ),
( 1763 ),
( 1766 ),
( 1769 ),
( 1772 ),
( 1775 ),
( 1778 ),
( 1781 ),
( 1784 ),
( 1787 ),
( 1790 ),
( 1793 ),
( 1795 ),
( 1798 ),
( 1801 ),
( 1804 ),
( 1807 ),
( 1810 ),
( 1813 ),
( 1817 ),
( 1820 ),
( 1823 ),
( 1826 ),
( 1829 ),
( 1832 ),
( 1835 ),
( 1838 ),
( 1841 ),
( 1844 ),
( 1847 ),
( 1851 ),
( 1854 ),
( 1857 ),
( 1860 ),
( 1863 ),
( 1867 ),
( 1870 ),
( 1873 ),
( 1876 ),
( 1879 ),
( 1883 ),
( 1886 ),
( 1889 ),
( 1893 ),
( 1896 ),
( 1899 ),
( 1903 ),
( 1906 ),
( 1909 ),
( 1913 ),
( 1916 ),
( 1919 ),
( 1923 ),
( 1926 ),
( 1930 ),
( 1933 ),
( 1936 ),
( 1940 ),
( 1943 ),
( 1947 ),
( 1950 ),
( 1954 ),
( 1957 ),
( 1961 ),
( 1965 ),
( 1968 ),
( 1972 ),
( 1975 ),
( 1979 ),
( 1982 ),
( 1986 ),
( 1990 ),
( 1993 ),
( 1997 ),
( 2001 ),
( 2004 ),
( 2008 ),
( 2012 ),
( 2016 ),
( 2019 ),
( 2023 ),
( 2027 ),
( 2031 ),
( 2035 ),
( 2038 ),
( 2042 ),
( 2046 ),
( 2050 ),
( 2054 ),
( 2058 ),
( 2062 ),
( 2065 ),
( 2069 ),
( 2073 ),
( 2077 ),
( 2081 ),
( 2085 ),
( 2089 ),
( 2093 ),
( 2097 ),
( 2101 ),
( 2106 ),
( 2110 ),
( 2114 ),
( 2118 ),
( 2122 ),
( 2126 ),
( 2130 ),
( 2135 ),
( 2139 ),
( 2143 ),
( 2147 ),
( 2151 ),
( 2156 ),
( 2160 ),
( 2164 ),
( 2169 ),
( 2173 ),
( 2177 ),
( 2182 ),
( 2186 ),
( 2191 ),
( 2195 ),
( 2199 ),
( 2204 ),
( 2208 ),
( 2213 ),
( 2217 ),
( 2222 ),
( 2227 ),
( 2231 ),
( 2236 ),
( 2240 ),
( 2245 ),
( 2250 ),
( 2254 ),
( 2259 ),
( 2264 ),
( 2268 ),
( 2273 ),
( 2278 ),
( 2283 ),
( 2288 ),
( 2292 ),
( 2297 ),
( 2302 ),
( 2307 ),
( 2312 ),
( 2317 ),
( 2322 ),
( 2327 ),
( 2332 ),
( 2337 ),
( 2342 ),
( 2347 ),
( 2352 ),
( 2357 ),
( 2362 ),
( 2367 ),
( 2373 ),
( 2378 ),
( 2383 ),
( 2388 ),
( 2394 ),
( 2399 ),
( 2404 ),
( 2409 ),
( 2415 ),
( 2420 ),
( 2426 ),
( 2431 ),
( 2437 ),
( 2442 ),
( 2448 ),
( 2453 ),
( 2459 ),
( 2464 ),
( 2470 ),
( 2475 ),
( 2481 ),
( 2487 ),
( 2493 ),
( 2498 ),
( 2504 ),
( 2510 ),
( 2516 ),
( 2521 ),
( 2527 ),
( 2533 ),
( 2539 ),
( 2545 ),
( 2551 ),
( 2557 ),
( 2563 ),
( 2569 ),
( 2575 ),
( 2581 ),
( 2588 ),
( 2594 ),
( 2600 ),
( 2606 ),
( 2613 ),
( 2619 ),
( 2625 ),
( 2632 ),
( 2638 ),
( 2644 ),
( 2651 ),
( 2657 ),
( 2664 ),
( 2670 ),
( 2677 ),
( 2684 ),
( 2690 ),
( 2697 ),
( 2704 ),
( 2710 ),
( 2717 ),
( 2724 ),
( 2731 ),
( 2738 ),
( 2745 ),
( 2752 ),
( 2759 ),
( 2766 ),
( 2773 ),
( 2780 ),
( 2787 ),
( 2794 ),
( 2801 ),
( 2809 ),
( 2816 ),
( 2823 ),
( 2831 ),
( 2838 ),
( 2845 ),
( 2853 ),
( 2860 ),
( 2868 ),
( 2876 ),
( 2883 ),
( 2891 ),
( 2899 ),
( 2906 ),
( 2914 ),
( 2922 ),
( 2930 ),
( 2938 ),
( 2946 ),
( 2954 ),
( 2962 ),
( 2970 ),
( 2978 ),
( 2986 ),
( 2995 ),
( 3003 ),
( 3011 ),
( 3020 ),
( 3028 ),
( 3037 ),
( 3045 ),
( 3054 ),
( 3062 ),
( 3071 ),
( 3080 ),
( 3088 ),
( 3097 ),
( 3106 ),
( 3115 ),
( 3124 ),
( 3133 ),
( 3142 ),
( 3151 ),
( 3160 ),
( 3170 ),
( 3179 ),
( 3188 ),
( 3198 ),
( 3207 ),
( 3217 ),
( 3226 ),
( 3236 ),
( 3245 ),
( 3255 ),
( 3265 ),
( 3275 ),
( 3285 ),
( 3295 ),
( 3305 ),
( 3315 ),
( 3325 ),
( 3335 ),
( 3346 ),
( 3356 ),
( 3366 ),
( 3377 ),
( 3387 ),
( 3398 ),
( 3409 ),
( 3419 ),
( 3430 ),
( 3441 ),
( 3452 ),
( 3463 ),
( 3474 ),
( 3485 ),
( 3496 ),
( 3508 ),
( 3519 ),
( 3531 ),
( 3542 ),
( 3554 ),
( 3565 ),
( 3577 ),
( 3589 ),
( 3601 ),
( 3613 ),
( 3625 ),
( 3637 ),
( 3649 ),
( 3662 ),
( 3674 ),
( 3687 ),
( 3699 ),
( 3712 ),
( 3724 ),
( 3737 ),
( 3750 ),
( 3763 ),
( 3776 ),
( 3790 ),
( 3803 ),
( 3816 ),
( 3830 ),
( 3843 ),
( 3857 ),
( 3871 ),
( 3884 ),
( 3898 ),
( 3913 ),
( 3927 ),
( 3941 ),
( 3955 ),
( 3970 ),
( 3984 ),
( 3999 ),
( 4014 ),
( 4029 ),
( 4044 ),
( 4059 ),
( 4074 ),
( 4089 ),
( 4105 ),
( 4121 ),
( 4136 ),
( 4152 ),
( 4168 ),
( 4184 ),
( 4200 ),
( 4217 ),
( 4233 ),
( 4250 ),
( 4266 ),
( 4283 ),
( 4300 ),
( 4317 ),
( 4334 ),
( 4352 ),
( 4369 ),
( 4387 ),
( 4405 ),
( 4423 ),
( 4441 ),
( 4459 ),
( 4478 ),
( 4496 ),
( 4515 ),
( 4534 ),
( 4553 ),
( 4572 ),
( 4591 ),
( 4611 ),
( 4630 ),
( 4650 ),
( 4670 ),
( 4691 ),
( 4711 ),
( 4731 ),
( 4752 ),
( 4773 ),
( 4794 ),
( 4815 ),
( 4837 ),
( 4859 ),
( 4880 ),
( 4902 ),
( 4925 ),
( 4947 ),
( 4970 ),
( 4993 ),
( 5016 ),
( 5039 ),
( 5063 ),
( 5086 ),
( 5110 ),
( 5134 ),
( 5159 ),
( 5183 ),
( 5208 ),
( 5233 ),
( 5259 ),
( 5284 ),
( 5310 ),
( 5336 ),
( 5363 ),
( 5389 ),
( 5416 ),
( 5443 ),
( 5471 ),
( 5499 ),
( 5527 ),
( 5555 ),
( 5584 ),
( 5612 ),
( 5642 ),
( 5671 ),
( 5701 ),
( 5731 ),
( 5761 ),
( 5792 ),
( 5823 ),
( 5855 ),
( 5886 ),
( 5919 ),
( 5951 ),
( 5984 ),
( 6017 ),
( 6051 ),
( 6085 ),
( 6119 ),
( 6154 ),
( 6189 ),
( 6224 ),
( 6260 ),
( 6296 ),
( 6333 ),
( 6370 ),
( 6408 ),
( 6446 ),
( 6484 ),
( 6523 ),
( 6563 ),
( 6603 ),
( 6643 ),
( 6684 ),
( 6726 ),
( 6768 ),
( 6810 ),
( 6853 ),
( 6897 ),
( 6941 ),
( 6985 ),
( 7031 ),
( 7077 ),
( 7123 ),
( 7170 ),
( 7218 ),
( 7266 ),
( 7315 ),
( 7365 ),
( 7415 ),
( 7466 ),
( 7518 ),
( 7570 ),
( 7623 ),
( 7677 ),
( 7732 ),
( 7788 ),
( 7844 ),
( 7901 ),
( 7959 ),
( 8018 ),
( 8077 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 ),
( 6103 )
);


--Eqn 50,000,000/ (4*(49700/9)-(47x/36))
--Where x is the distance ranging from 400 mm to 4000mm
-- x<=400mm then the period = 50,000,000/(4 * 5000Hz))  
-- x>=4000mm then the period = 50,000,000/(4 * 30Hz)) 
constant d2b_LUT : array_1d := (
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2500 ),
( 2501 ),
( 2501 ),
( 2502 ),
( 2503 ),
( 2503 ),
( 2504 ),
( 2505 ),
( 2505 ),
( 2506 ),
( 2507 ),
( 2507 ),
( 2508 ),
( 2509 ),
( 2509 ),
( 2510 ),
( 2511 ),
( 2511 ),
( 2512 ),
( 2513 ),
( 2513 ),
( 2514 ),
( 2515 ),
( 2515 ),
( 2516 ),
( 2517 ),
( 2517 ),
( 2518 ),
( 2519 ),
( 2519 ),
( 2520 ),
( 2521 ),
( 2521 ),
( 2522 ),
( 2523 ),
( 2523 ),
( 2524 ),
( 2525 ),
( 2525 ),
( 2526 ),
( 2527 ),
( 2527 ),
( 2528 ),
( 2529 ),
( 2529 ),
( 2530 ),
( 2531 ),
( 2531 ),
( 2532 ),
( 2533 ),
( 2533 ),
( 2534 ),
( 2535 ),
( 2535 ),
( 2536 ),
( 2537 ),
( 2537 ),
( 2538 ),
( 2539 ),
( 2539 ),
( 2540 ),
( 2541 ),
( 2541 ),
( 2542 ),
( 2543 ),
( 2543 ),
( 2544 ),
( 2545 ),
( 2545 ),
( 2546 ),
( 2547 ),
( 2547 ),
( 2548 ),
( 2549 ),
( 2549 ),
( 2550 ),
( 2551 ),
( 2551 ),
( 2552 ),
( 2553 ),
( 2553 ),
( 2554 ),
( 2555 ),
( 2555 ),
( 2556 ),
( 2557 ),
( 2558 ),
( 2558 ),
( 2559 ),
( 2560 ),
( 2560 ),
( 2561 ),
( 2562 ),
( 2562 ),
( 2563 ),
( 2564 ),
( 2564 ),
( 2565 ),
( 2566 ),
( 2566 ),
( 2567 ),
( 2568 ),
( 2569 ),
( 2569 ),
( 2570 ),
( 2571 ),
( 2571 ),
( 2572 ),
( 2573 ),
( 2573 ),
( 2574 ),
( 2575 ),
( 2575 ),
( 2576 ),
( 2577 ),
( 2578 ),
( 2578 ),
( 2579 ),
( 2580 ),
( 2580 ),
( 2581 ),
( 2582 ),
( 2582 ),
( 2583 ),
( 2584 ),
( 2584 ),
( 2585 ),
( 2586 ),
( 2587 ),
( 2587 ),
( 2588 ),
( 2589 ),
( 2589 ),
( 2590 ),
( 2591 ),
( 2591 ),
( 2592 ),
( 2593 ),
( 2594 ),
( 2594 ),
( 2595 ),
( 2596 ),
( 2596 ),
( 2597 ),
( 2598 ),
( 2598 ),
( 2599 ),
( 2600 ),
( 2601 ),
( 2601 ),
( 2602 ),
( 2603 ),
( 2603 ),
( 2604 ),
( 2605 ),
( 2606 ),
( 2606 ),
( 2607 ),
( 2608 ),
( 2608 ),
( 2609 ),
( 2610 ),
( 2611 ),
( 2611 ),
( 2612 ),
( 2613 ),
( 2613 ),
( 2614 ),
( 2615 ),
( 2616 ),
( 2616 ),
( 2617 ),
( 2618 ),
( 2618 ),
( 2619 ),
( 2620 ),
( 2621 ),
( 2621 ),
( 2622 ),
( 2623 ),
( 2623 ),
( 2624 ),
( 2625 ),
( 2626 ),
( 2626 ),
( 2627 ),
( 2628 ),
( 2628 ),
( 2629 ),
( 2630 ),
( 2631 ),
( 2631 ),
( 2632 ),
( 2633 ),
( 2634 ),
( 2634 ),
( 2635 ),
( 2636 ),
( 2636 ),
( 2637 ),
( 2638 ),
( 2639 ),
( 2639 ),
( 2640 ),
( 2641 ),
( 2642 ),
( 2642 ),
( 2643 ),
( 2644 ),
( 2644 ),
( 2645 ),
( 2646 ),
( 2647 ),
( 2647 ),
( 2648 ),
( 2649 ),
( 2650 ),
( 2650 ),
( 2651 ),
( 2652 ),
( 2652 ),
( 2653 ),
( 2654 ),
( 2655 ),
( 2655 ),
( 2656 ),
( 2657 ),
( 2658 ),
( 2658 ),
( 2659 ),
( 2660 ),
( 2661 ),
( 2661 ),
( 2662 ),
( 2663 ),
( 2664 ),
( 2664 ),
( 2665 ),
( 2666 ),
( 2667 ),
( 2667 ),
( 2668 ),
( 2669 ),
( 2669 ),
( 2670 ),
( 2671 ),
( 2672 ),
( 2672 ),
( 2673 ),
( 2674 ),
( 2675 ),
( 2675 ),
( 2676 ),
( 2677 ),
( 2678 ),
( 2678 ),
( 2679 ),
( 2680 ),
( 2681 ),
( 2681 ),
( 2682 ),
( 2683 ),
( 2684 ),
( 2684 ),
( 2685 ),
( 2686 ),
( 2687 ),
( 2687 ),
( 2688 ),
( 2689 ),
( 2690 ),
( 2691 ),
( 2691 ),
( 2692 ),
( 2693 ),
( 2694 ),
( 2694 ),
( 2695 ),
( 2696 ),
( 2697 ),
( 2697 ),
( 2698 ),
( 2699 ),
( 2700 ),
( 2700 ),
( 2701 ),
( 2702 ),
( 2703 ),
( 2703 ),
( 2704 ),
( 2705 ),
( 2706 ),
( 2706 ),
( 2707 ),
( 2708 ),
( 2709 ),
( 2710 ),
( 2710 ),
( 2711 ),
( 2712 ),
( 2713 ),
( 2713 ),
( 2714 ),
( 2715 ),
( 2716 ),
( 2716 ),
( 2717 ),
( 2718 ),
( 2719 ),
( 2720 ),
( 2720 ),
( 2721 ),
( 2722 ),
( 2723 ),
( 2723 ),
( 2724 ),
( 2725 ),
( 2726 ),
( 2727 ),
( 2727 ),
( 2728 ),
( 2729 ),
( 2730 ),
( 2730 ),
( 2731 ),
( 2732 ),
( 2733 ),
( 2734 ),
( 2734 ),
( 2735 ),
( 2736 ),
( 2737 ),
( 2737 ),
( 2738 ),
( 2739 ),
( 2740 ),
( 2741 ),
( 2741 ),
( 2742 ),
( 2743 ),
( 2744 ),
( 2744 ),
( 2745 ),
( 2746 ),
( 2747 ),
( 2748 ),
( 2748 ),
( 2749 ),
( 2750 ),
( 2751 ),
( 2752 ),
( 2752 ),
( 2753 ),
( 2754 ),
( 2755 ),
( 2756 ),
( 2756 ),
( 2757 ),
( 2758 ),
( 2759 ),
( 2760 ),
( 2760 ),
( 2761 ),
( 2762 ),
( 2763 ),
( 2763 ),
( 2764 ),
( 2765 ),
( 2766 ),
( 2767 ),
( 2767 ),
( 2768 ),
( 2769 ),
( 2770 ),
( 2771 ),
( 2771 ),
( 2772 ),
( 2773 ),
( 2774 ),
( 2775 ),
( 2776 ),
( 2776 ),
( 2777 ),
( 2778 ),
( 2779 ),
( 2780 ),
( 2780 ),
( 2781 ),
( 2782 ),
( 2783 ),
( 2784 ),
( 2784 ),
( 2785 ),
( 2786 ),
( 2787 ),
( 2788 ),
( 2788 ),
( 2789 ),
( 2790 ),
( 2791 ),
( 2792 ),
( 2793 ),
( 2793 ),
( 2794 ),
( 2795 ),
( 2796 ),
( 2797 ),
( 2797 ),
( 2798 ),
( 2799 ),
( 2800 ),
( 2801 ),
( 2802 ),
( 2802 ),
( 2803 ),
( 2804 ),
( 2805 ),
( 2806 ),
( 2806 ),
( 2807 ),
( 2808 ),
( 2809 ),
( 2810 ),
( 2811 ),
( 2811 ),
( 2812 ),
( 2813 ),
( 2814 ),
( 2815 ),
( 2816 ),
( 2816 ),
( 2817 ),
( 2818 ),
( 2819 ),
( 2820 ),
( 2820 ),
( 2821 ),
( 2822 ),
( 2823 ),
( 2824 ),
( 2825 ),
( 2825 ),
( 2826 ),
( 2827 ),
( 2828 ),
( 2829 ),
( 2830 ),
( 2830 ),
( 2831 ),
( 2832 ),
( 2833 ),
( 2834 ),
( 2835 ),
( 2836 ),
( 2836 ),
( 2837 ),
( 2838 ),
( 2839 ),
( 2840 ),
( 2841 ),
( 2841 ),
( 2842 ),
( 2843 ),
( 2844 ),
( 2845 ),
( 2846 ),
( 2846 ),
( 2847 ),
( 2848 ),
( 2849 ),
( 2850 ),
( 2851 ),
( 2852 ),
( 2852 ),
( 2853 ),
( 2854 ),
( 2855 ),
( 2856 ),
( 2857 ),
( 2858 ),
( 2858 ),
( 2859 ),
( 2860 ),
( 2861 ),
( 2862 ),
( 2863 ),
( 2864 ),
( 2864 ),
( 2865 ),
( 2866 ),
( 2867 ),
( 2868 ),
( 2869 ),
( 2870 ),
( 2870 ),
( 2871 ),
( 2872 ),
( 2873 ),
( 2874 ),
( 2875 ),
( 2876 ),
( 2876 ),
( 2877 ),
( 2878 ),
( 2879 ),
( 2880 ),
( 2881 ),
( 2882 ),
( 2882 ),
( 2883 ),
( 2884 ),
( 2885 ),
( 2886 ),
( 2887 ),
( 2888 ),
( 2889 ),
( 2889 ),
( 2890 ),
( 2891 ),
( 2892 ),
( 2893 ),
( 2894 ),
( 2895 ),
( 2896 ),
( 2896 ),
( 2897 ),
( 2898 ),
( 2899 ),
( 2900 ),
( 2901 ),
( 2902 ),
( 2903 ),
( 2903 ),
( 2904 ),
( 2905 ),
( 2906 ),
( 2907 ),
( 2908 ),
( 2909 ),
( 2910 ),
( 2911 ),
( 2911 ),
( 2912 ),
( 2913 ),
( 2914 ),
( 2915 ),
( 2916 ),
( 2917 ),
( 2918 ),
( 2918 ),
( 2919 ),
( 2920 ),
( 2921 ),
( 2922 ),
( 2923 ),
( 2924 ),
( 2925 ),
( 2926 ),
( 2927 ),
( 2927 ),
( 2928 ),
( 2929 ),
( 2930 ),
( 2931 ),
( 2932 ),
( 2933 ),
( 2934 ),
( 2935 ),
( 2935 ),
( 2936 ),
( 2937 ),
( 2938 ),
( 2939 ),
( 2940 ),
( 2941 ),
( 2942 ),
( 2943 ),
( 2944 ),
( 2945 ),
( 2945 ),
( 2946 ),
( 2947 ),
( 2948 ),
( 2949 ),
( 2950 ),
( 2951 ),
( 2952 ),
( 2953 ),
( 2954 ),
( 2955 ),
( 2955 ),
( 2956 ),
( 2957 ),
( 2958 ),
( 2959 ),
( 2960 ),
( 2961 ),
( 2962 ),
( 2963 ),
( 2964 ),
( 2965 ),
( 2966 ),
( 2966 ),
( 2967 ),
( 2968 ),
( 2969 ),
( 2970 ),
( 2971 ),
( 2972 ),
( 2973 ),
( 2974 ),
( 2975 ),
( 2976 ),
( 2977 ),
( 2977 ),
( 2978 ),
( 2979 ),
( 2980 ),
( 2981 ),
( 2982 ),
( 2983 ),
( 2984 ),
( 2985 ),
( 2986 ),
( 2987 ),
( 2988 ),
( 2989 ),
( 2990 ),
( 2991 ),
( 2991 ),
( 2992 ),
( 2993 ),
( 2994 ),
( 2995 ),
( 2996 ),
( 2997 ),
( 2998 ),
( 2999 ),
( 3000 ),
( 3001 ),
( 3002 ),
( 3003 ),
( 3004 ),
( 3005 ),
( 3006 ),
( 3006 ),
( 3007 ),
( 3008 ),
( 3009 ),
( 3010 ),
( 3011 ),
( 3012 ),
( 3013 ),
( 3014 ),
( 3015 ),
( 3016 ),
( 3017 ),
( 3018 ),
( 3019 ),
( 3020 ),
( 3021 ),
( 3022 ),
( 3023 ),
( 3024 ),
( 3025 ),
( 3025 ),
( 3026 ),
( 3027 ),
( 3028 ),
( 3029 ),
( 3030 ),
( 3031 ),
( 3032 ),
( 3033 ),
( 3034 ),
( 3035 ),
( 3036 ),
( 3037 ),
( 3038 ),
( 3039 ),
( 3040 ),
( 3041 ),
( 3042 ),
( 3043 ),
( 3044 ),
( 3045 ),
( 3046 ),
( 3047 ),
( 3048 ),
( 3049 ),
( 3050 ),
( 3051 ),
( 3052 ),
( 3052 ),
( 3053 ),
( 3054 ),
( 3055 ),
( 3056 ),
( 3057 ),
( 3058 ),
( 3059 ),
( 3060 ),
( 3061 ),
( 3062 ),
( 3063 ),
( 3064 ),
( 3065 ),
( 3066 ),
( 3067 ),
( 3068 ),
( 3069 ),
( 3070 ),
( 3071 ),
( 3072 ),
( 3073 ),
( 3074 ),
( 3075 ),
( 3076 ),
( 3077 ),
( 3078 ),
( 3079 ),
( 3080 ),
( 3081 ),
( 3082 ),
( 3083 ),
( 3084 ),
( 3085 ),
( 3086 ),
( 3087 ),
( 3088 ),
( 3089 ),
( 3090 ),
( 3091 ),
( 3092 ),
( 3093 ),
( 3094 ),
( 3095 ),
( 3096 ),
( 3097 ),
( 3098 ),
( 3099 ),
( 3100 ),
( 3101 ),
( 3102 ),
( 3103 ),
( 3104 ),
( 3105 ),
( 3106 ),
( 3107 ),
( 3108 ),
( 3109 ),
( 3110 ),
( 3111 ),
( 3112 ),
( 3113 ),
( 3114 ),
( 3115 ),
( 3116 ),
( 3117 ),
( 3118 ),
( 3119 ),
( 3120 ),
( 3121 ),
( 3122 ),
( 3123 ),
( 3124 ),
( 3125 ),
( 3126 ),
( 3127 ),
( 3128 ),
( 3129 ),
( 3130 ),
( 3131 ),
( 3132 ),
( 3133 ),
( 3134 ),
( 3135 ),
( 3136 ),
( 3138 ),
( 3139 ),
( 3140 ),
( 3141 ),
( 3142 ),
( 3143 ),
( 3144 ),
( 3145 ),
( 3146 ),
( 3147 ),
( 3148 ),
( 3149 ),
( 3150 ),
( 3151 ),
( 3152 ),
( 3153 ),
( 3154 ),
( 3155 ),
( 3156 ),
( 3157 ),
( 3158 ),
( 3159 ),
( 3160 ),
( 3161 ),
( 3162 ),
( 3163 ),
( 3164 ),
( 3166 ),
( 3167 ),
( 3168 ),
( 3169 ),
( 3170 ),
( 3171 ),
( 3172 ),
( 3173 ),
( 3174 ),
( 3175 ),
( 3176 ),
( 3177 ),
( 3178 ),
( 3179 ),
( 3180 ),
( 3181 ),
( 3182 ),
( 3183 ),
( 3184 ),
( 3186 ),
( 3187 ),
( 3188 ),
( 3189 ),
( 3190 ),
( 3191 ),
( 3192 ),
( 3193 ),
( 3194 ),
( 3195 ),
( 3196 ),
( 3197 ),
( 3198 ),
( 3199 ),
( 3200 ),
( 3202 ),
( 3203 ),
( 3204 ),
( 3205 ),
( 3206 ),
( 3207 ),
( 3208 ),
( 3209 ),
( 3210 ),
( 3211 ),
( 3212 ),
( 3213 ),
( 3214 ),
( 3215 ),
( 3217 ),
( 3218 ),
( 3219 ),
( 3220 ),
( 3221 ),
( 3222 ),
( 3223 ),
( 3224 ),
( 3225 ),
( 3226 ),
( 3227 ),
( 3228 ),
( 3230 ),
( 3231 ),
( 3232 ),
( 3233 ),
( 3234 ),
( 3235 ),
( 3236 ),
( 3237 ),
( 3238 ),
( 3239 ),
( 3241 ),
( 3242 ),
( 3243 ),
( 3244 ),
( 3245 ),
( 3246 ),
( 3247 ),
( 3248 ),
( 3249 ),
( 3250 ),
( 3252 ),
( 3253 ),
( 3254 ),
( 3255 ),
( 3256 ),
( 3257 ),
( 3258 ),
( 3259 ),
( 3260 ),
( 3261 ),
( 3263 ),
( 3264 ),
( 3265 ),
( 3266 ),
( 3267 ),
( 3268 ),
( 3269 ),
( 3270 ),
( 3272 ),
( 3273 ),
( 3274 ),
( 3275 ),
( 3276 ),
( 3277 ),
( 3278 ),
( 3279 ),
( 3280 ),
( 3282 ),
( 3283 ),
( 3284 ),
( 3285 ),
( 3286 ),
( 3287 ),
( 3288 ),
( 3289 ),
( 3291 ),
( 3292 ),
( 3293 ),
( 3294 ),
( 3295 ),
( 3296 ),
( 3297 ),
( 3299 ),
( 3300 ),
( 3301 ),
( 3302 ),
( 3303 ),
( 3304 ),
( 3305 ),
( 3307 ),
( 3308 ),
( 3309 ),
( 3310 ),
( 3311 ),
( 3312 ),
( 3313 ),
( 3315 ),
( 3316 ),
( 3317 ),
( 3318 ),
( 3319 ),
( 3320 ),
( 3321 ),
( 3323 ),
( 3324 ),
( 3325 ),
( 3326 ),
( 3327 ),
( 3328 ),
( 3330 ),
( 3331 ),
( 3332 ),
( 3333 ),
( 3334 ),
( 3335 ),
( 3336 ),
( 3338 ),
( 3339 ),
( 3340 ),
( 3341 ),
( 3342 ),
( 3343 ),
( 3345 ),
( 3346 ),
( 3347 ),
( 3348 ),
( 3349 ),
( 3351 ),
( 3352 ),
( 3353 ),
( 3354 ),
( 3355 ),
( 3356 ),
( 3358 ),
( 3359 ),
( 3360 ),
( 3361 ),
( 3362 ),
( 3363 ),
( 3365 ),
( 3366 ),
( 3367 ),
( 3368 ),
( 3369 ),
( 3371 ),
( 3372 ),
( 3373 ),
( 3374 ),
( 3375 ),
( 3377 ),
( 3378 ),
( 3379 ),
( 3380 ),
( 3381 ),
( 3382 ),
( 3384 ),
( 3385 ),
( 3386 ),
( 3387 ),
( 3388 ),
( 3390 ),
( 3391 ),
( 3392 ),
( 3393 ),
( 3394 ),
( 3396 ),
( 3397 ),
( 3398 ),
( 3399 ),
( 3400 ),
( 3402 ),
( 3403 ),
( 3404 ),
( 3405 ),
( 3407 ),
( 3408 ),
( 3409 ),
( 3410 ),
( 3411 ),
( 3413 ),
( 3414 ),
( 3415 ),
( 3416 ),
( 3417 ),
( 3419 ),
( 3420 ),
( 3421 ),
( 3422 ),
( 3424 ),
( 3425 ),
( 3426 ),
( 3427 ),
( 3428 ),
( 3430 ),
( 3431 ),
( 3432 ),
( 3433 ),
( 3435 ),
( 3436 ),
( 3437 ),
( 3438 ),
( 3440 ),
( 3441 ),
( 3442 ),
( 3443 ),
( 3445 ),
( 3446 ),
( 3447 ),
( 3448 ),
( 3449 ),
( 3451 ),
( 3452 ),
( 3453 ),
( 3454 ),
( 3456 ),
( 3457 ),
( 3458 ),
( 3459 ),
( 3461 ),
( 3462 ),
( 3463 ),
( 3464 ),
( 3466 ),
( 3467 ),
( 3468 ),
( 3469 ),
( 3471 ),
( 3472 ),
( 3473 ),
( 3475 ),
( 3476 ),
( 3477 ),
( 3478 ),
( 3480 ),
( 3481 ),
( 3482 ),
( 3483 ),
( 3485 ),
( 3486 ),
( 3487 ),
( 3488 ),
( 3490 ),
( 3491 ),
( 3492 ),
( 3494 ),
( 3495 ),
( 3496 ),
( 3497 ),
( 3499 ),
( 3500 ),
( 3501 ),
( 3502 ),
( 3504 ),
( 3505 ),
( 3506 ),
( 3508 ),
( 3509 ),
( 3510 ),
( 3511 ),
( 3513 ),
( 3514 ),
( 3515 ),
( 3517 ),
( 3518 ),
( 3519 ),
( 3521 ),
( 3522 ),
( 3523 ),
( 3524 ),
( 3526 ),
( 3527 ),
( 3528 ),
( 3530 ),
( 3531 ),
( 3532 ),
( 3534 ),
( 3535 ),
( 3536 ),
( 3537 ),
( 3539 ),
( 3540 ),
( 3541 ),
( 3543 ),
( 3544 ),
( 3545 ),
( 3547 ),
( 3548 ),
( 3549 ),
( 3551 ),
( 3552 ),
( 3553 ),
( 3555 ),
( 3556 ),
( 3557 ),
( 3558 ),
( 3560 ),
( 3561 ),
( 3562 ),
( 3564 ),
( 3565 ),
( 3566 ),
( 3568 ),
( 3569 ),
( 3570 ),
( 3572 ),
( 3573 ),
( 3574 ),
( 3576 ),
( 3577 ),
( 3578 ),
( 3580 ),
( 3581 ),
( 3582 ),
( 3584 ),
( 3585 ),
( 3586 ),
( 3588 ),
( 3589 ),
( 3590 ),
( 3592 ),
( 3593 ),
( 3595 ),
( 3596 ),
( 3597 ),
( 3599 ),
( 3600 ),
( 3601 ),
( 3603 ),
( 3604 ),
( 3605 ),
( 3607 ),
( 3608 ),
( 3609 ),
( 3611 ),
( 3612 ),
( 3614 ),
( 3615 ),
( 3616 ),
( 3618 ),
( 3619 ),
( 3620 ),
( 3622 ),
( 3623 ),
( 3624 ),
( 3626 ),
( 3627 ),
( 3629 ),
( 3630 ),
( 3631 ),
( 3633 ),
( 3634 ),
( 3635 ),
( 3637 ),
( 3638 ),
( 3640 ),
( 3641 ),
( 3642 ),
( 3644 ),
( 3645 ),
( 3647 ),
( 3648 ),
( 3649 ),
( 3651 ),
( 3652 ),
( 3654 ),
( 3655 ),
( 3656 ),
( 3658 ),
( 3659 ),
( 3661 ),
( 3662 ),
( 3663 ),
( 3665 ),
( 3666 ),
( 3668 ),
( 3669 ),
( 3670 ),
( 3672 ),
( 3673 ),
( 3675 ),
( 3676 ),
( 3677 ),
( 3679 ),
( 3680 ),
( 3682 ),
( 3683 ),
( 3684 ),
( 3686 ),
( 3687 ),
( 3689 ),
( 3690 ),
( 3692 ),
( 3693 ),
( 3694 ),
( 3696 ),
( 3697 ),
( 3699 ),
( 3700 ),
( 3702 ),
( 3703 ),
( 3704 ),
( 3706 ),
( 3707 ),
( 3709 ),
( 3710 ),
( 3712 ),
( 3713 ),
( 3714 ),
( 3716 ),
( 3717 ),
( 3719 ),
( 3720 ),
( 3722 ),
( 3723 ),
( 3725 ),
( 3726 ),
( 3727 ),
( 3729 ),
( 3730 ),
( 3732 ),
( 3733 ),
( 3735 ),
( 3736 ),
( 3738 ),
( 3739 ),
( 3741 ),
( 3742 ),
( 3744 ),
( 3745 ),
( 3746 ),
( 3748 ),
( 3749 ),
( 3751 ),
( 3752 ),
( 3754 ),
( 3755 ),
( 3757 ),
( 3758 ),
( 3760 ),
( 3761 ),
( 3763 ),
( 3764 ),
( 3766 ),
( 3767 ),
( 3769 ),
( 3770 ),
( 3772 ),
( 3773 ),
( 3775 ),
( 3776 ),
( 3777 ),
( 3779 ),
( 3780 ),
( 3782 ),
( 3783 ),
( 3785 ),
( 3786 ),
( 3788 ),
( 3789 ),
( 3791 ),
( 3792 ),
( 3794 ),
( 3795 ),
( 3797 ),
( 3798 ),
( 3800 ),
( 3801 ),
( 3803 ),
( 3804 ),
( 3806 ),
( 3808 ),
( 3809 ),
( 3811 ),
( 3812 ),
( 3814 ),
( 3815 ),
( 3817 ),
( 3818 ),
( 3820 ),
( 3821 ),
( 3823 ),
( 3824 ),
( 3826 ),
( 3827 ),
( 3829 ),
( 3830 ),
( 3832 ),
( 3833 ),
( 3835 ),
( 3837 ),
( 3838 ),
( 3840 ),
( 3841 ),
( 3843 ),
( 3844 ),
( 3846 ),
( 3847 ),
( 3849 ),
( 3850 ),
( 3852 ),
( 3853 ),
( 3855 ),
( 3857 ),
( 3858 ),
( 3860 ),
( 3861 ),
( 3863 ),
( 3864 ),
( 3866 ),
( 3868 ),
( 3869 ),
( 3871 ),
( 3872 ),
( 3874 ),
( 3875 ),
( 3877 ),
( 3878 ),
( 3880 ),
( 3882 ),
( 3883 ),
( 3885 ),
( 3886 ),
( 3888 ),
( 3890 ),
( 3891 ),
( 3893 ),
( 3894 ),
( 3896 ),
( 3897 ),
( 3899 ),
( 3901 ),
( 3902 ),
( 3904 ),
( 3905 ),
( 3907 ),
( 3909 ),
( 3910 ),
( 3912 ),
( 3913 ),
( 3915 ),
( 3917 ),
( 3918 ),
( 3920 ),
( 3921 ),
( 3923 ),
( 3925 ),
( 3926 ),
( 3928 ),
( 3929 ),
( 3931 ),
( 3933 ),
( 3934 ),
( 3936 ),
( 3937 ),
( 3939 ),
( 3941 ),
( 3942 ),
( 3944 ),
( 3946 ),
( 3947 ),
( 3949 ),
( 3950 ),
( 3952 ),
( 3954 ),
( 3955 ),
( 3957 ),
( 3959 ),
( 3960 ),
( 3962 ),
( 3964 ),
( 3965 ),
( 3967 ),
( 3968 ),
( 3970 ),
( 3972 ),
( 3973 ),
( 3975 ),
( 3977 ),
( 3978 ),
( 3980 ),
( 3982 ),
( 3983 ),
( 3985 ),
( 3987 ),
( 3988 ),
( 3990 ),
( 3992 ),
( 3993 ),
( 3995 ),
( 3997 ),
( 3998 ),
( 4000 ),
( 4002 ),
( 4003 ),
( 4005 ),
( 4007 ),
( 4008 ),
( 4010 ),
( 4012 ),
( 4013 ),
( 4015 ),
( 4017 ),
( 4018 ),
( 4020 ),
( 4022 ),
( 4024 ),
( 4025 ),
( 4027 ),
( 4029 ),
( 4030 ),
( 4032 ),
( 4034 ),
( 4035 ),
( 4037 ),
( 4039 ),
( 4041 ),
( 4042 ),
( 4044 ),
( 4046 ),
( 4047 ),
( 4049 ),
( 4051 ),
( 4052 ),
( 4054 ),
( 4056 ),
( 4058 ),
( 4059 ),
( 4061 ),
( 4063 ),
( 4065 ),
( 4066 ),
( 4068 ),
( 4070 ),
( 4071 ),
( 4073 ),
( 4075 ),
( 4077 ),
( 4078 ),
( 4080 ),
( 4082 ),
( 4084 ),
( 4085 ),
( 4087 ),
( 4089 ),
( 4091 ),
( 4092 ),
( 4094 ),
( 4096 ),
( 4098 ),
( 4099 ),
( 4101 ),
( 4103 ),
( 4105 ),
( 4106 ),
( 4108 ),
( 4110 ),
( 4112 ),
( 4113 ),
( 4115 ),
( 4117 ),
( 4119 ),
( 4121 ),
( 4122 ),
( 4124 ),
( 4126 ),
( 4128 ),
( 4129 ),
( 4131 ),
( 4133 ),
( 4135 ),
( 4137 ),
( 4138 ),
( 4140 ),
( 4142 ),
( 4144 ),
( 4145 ),
( 4147 ),
( 4149 ),
( 4151 ),
( 4153 ),
( 4154 ),
( 4156 ),
( 4158 ),
( 4160 ),
( 4162 ),
( 4164 ),
( 4165 ),
( 4167 ),
( 4169 ),
( 4171 ),
( 4173 ),
( 4174 ),
( 4176 ),
( 4178 ),
( 4180 ),
( 4182 ),
( 4184 ),
( 4185 ),
( 4187 ),
( 4189 ),
( 4191 ),
( 4193 ),
( 4195 ),
( 4196 ),
( 4198 ),
( 4200 ),
( 4202 ),
( 4204 ),
( 4206 ),
( 4207 ),
( 4209 ),
( 4211 ),
( 4213 ),
( 4215 ),
( 4217 ),
( 4219 ),
( 4220 ),
( 4222 ),
( 4224 ),
( 4226 ),
( 4228 ),
( 4230 ),
( 4232 ),
( 4233 ),
( 4235 ),
( 4237 ),
( 4239 ),
( 4241 ),
( 4243 ),
( 4245 ),
( 4247 ),
( 4248 ),
( 4250 ),
( 4252 ),
( 4254 ),
( 4256 ),
( 4258 ),
( 4260 ),
( 4262 ),
( 4264 ),
( 4266 ),
( 4267 ),
( 4269 ),
( 4271 ),
( 4273 ),
( 4275 ),
( 4277 ),
( 4279 ),
( 4281 ),
( 4283 ),
( 4285 ),
( 4287 ),
( 4288 ),
( 4290 ),
( 4292 ),
( 4294 ),
( 4296 ),
( 4298 ),
( 4300 ),
( 4302 ),
( 4304 ),
( 4306 ),
( 4308 ),
( 4310 ),
( 4312 ),
( 4314 ),
( 4316 ),
( 4317 ),
( 4319 ),
( 4321 ),
( 4323 ),
( 4325 ),
( 4327 ),
( 4329 ),
( 4331 ),
( 4333 ),
( 4335 ),
( 4337 ),
( 4339 ),
( 4341 ),
( 4343 ),
( 4345 ),
( 4347 ),
( 4349 ),
( 4351 ),
( 4353 ),
( 4355 ),
( 4357 ),
( 4359 ),
( 4361 ),
( 4363 ),
( 4365 ),
( 4367 ),
( 4369 ),
( 4371 ),
( 4373 ),
( 4375 ),
( 4377 ),
( 4379 ),
( 4381 ),
( 4383 ),
( 4385 ),
( 4387 ),
( 4389 ),
( 4391 ),
( 4393 ),
( 4395 ),
( 4397 ),
( 4399 ),
( 4401 ),
( 4403 ),
( 4405 ),
( 4407 ),
( 4409 ),
( 4411 ),
( 4413 ),
( 4415 ),
( 4417 ),
( 4419 ),
( 4421 ),
( 4423 ),
( 4425 ),
( 4427 ),
( 4429 ),
( 4431 ),
( 4433 ),
( 4435 ),
( 4438 ),
( 4440 ),
( 4442 ),
( 4444 ),
( 4446 ),
( 4448 ),
( 4450 ),
( 4452 ),
( 4454 ),
( 4456 ),
( 4458 ),
( 4460 ),
( 4462 ),
( 4464 ),
( 4467 ),
( 4469 ),
( 4471 ),
( 4473 ),
( 4475 ),
( 4477 ),
( 4479 ),
( 4481 ),
( 4483 ),
( 4485 ),
( 4487 ),
( 4490 ),
( 4492 ),
( 4494 ),
( 4496 ),
( 4498 ),
( 4500 ),
( 4502 ),
( 4504 ),
( 4506 ),
( 4509 ),
( 4511 ),
( 4513 ),
( 4515 ),
( 4517 ),
( 4519 ),
( 4521 ),
( 4523 ),
( 4526 ),
( 4528 ),
( 4530 ),
( 4532 ),
( 4534 ),
( 4536 ),
( 4538 ),
( 4541 ),
( 4543 ),
( 4545 ),
( 4547 ),
( 4549 ),
( 4551 ),
( 4554 ),
( 4556 ),
( 4558 ),
( 4560 ),
( 4562 ),
( 4564 ),
( 4567 ),
( 4569 ),
( 4571 ),
( 4573 ),
( 4575 ),
( 4578 ),
( 4580 ),
( 4582 ),
( 4584 ),
( 4586 ),
( 4589 ),
( 4591 ),
( 4593 ),
( 4595 ),
( 4597 ),
( 4600 ),
( 4602 ),
( 4604 ),
( 4606 ),
( 4608 ),
( 4611 ),
( 4613 ),
( 4615 ),
( 4617 ),
( 4620 ),
( 4622 ),
( 4624 ),
( 4626 ),
( 4628 ),
( 4631 ),
( 4633 ),
( 4635 ),
( 4637 ),
( 4640 ),
( 4642 ),
( 4644 ),
( 4646 ),
( 4649 ),
( 4651 ),
( 4653 ),
( 4655 ),
( 4658 ),
( 4660 ),
( 4662 ),
( 4665 ),
( 4667 ),
( 4669 ),
( 4671 ),
( 4674 ),
( 4676 ),
( 4678 ),
( 4680 ),
( 4683 ),
( 4685 ),
( 4687 ),
( 4690 ),
( 4692 ),
( 4694 ),
( 4697 ),
( 4699 ),
( 4701 ),
( 4703 ),
( 4706 ),
( 4708 ),
( 4710 ),
( 4713 ),
( 4715 ),
( 4717 ),
( 4720 ),
( 4722 ),
( 4724 ),
( 4727 ),
( 4729 ),
( 4731 ),
( 4734 ),
( 4736 ),
( 4738 ),
( 4741 ),
( 4743 ),
( 4745 ),
( 4748 ),
( 4750 ),
( 4753 ),
( 4755 ),
( 4757 ),
( 4760 ),
( 4762 ),
( 4764 ),
( 4767 ),
( 4769 ),
( 4771 ),
( 4774 ),
( 4776 ),
( 4779 ),
( 4781 ),
( 4783 ),
( 4786 ),
( 4788 ),
( 4791 ),
( 4793 ),
( 4795 ),
( 4798 ),
( 4800 ),
( 4803 ),
( 4805 ),
( 4807 ),
( 4810 ),
( 4812 ),
( 4815 ),
( 4817 ),
( 4819 ),
( 4822 ),
( 4824 ),
( 4827 ),
( 4829 ),
( 4832 ),
( 4834 ),
( 4837 ),
( 4839 ),
( 4841 ),
( 4844 ),
( 4846 ),
( 4849 ),
( 4851 ),
( 4854 ),
( 4856 ),
( 4859 ),
( 4861 ),
( 4864 ),
( 4866 ),
( 4868 ),
( 4871 ),
( 4873 ),
( 4876 ),
( 4878 ),
( 4881 ),
( 4883 ),
( 4886 ),
( 4888 ),
( 4891 ),
( 4893 ),
( 4896 ),
( 4898 ),
( 4901 ),
( 4903 ),
( 4906 ),
( 4908 ),
( 4911 ),
( 4913 ),
( 4916 ),
( 4919 ),
( 4921 ),
( 4924 ),
( 4926 ),
( 4929 ),
( 4931 ),
( 4934 ),
( 4936 ),
( 4939 ),
( 4941 ),
( 4944 ),
( 4946 ),
( 4949 ),
( 4952 ),
( 4954 ),
( 4957 ),
( 4959 ),
( 4962 ),
( 4964 ),
( 4967 ),
( 4970 ),
( 4972 ),
( 4975 ),
( 4977 ),
( 4980 ),
( 4983 ),
( 4985 ),
( 4988 ),
( 4990 ),
( 4993 ),
( 4996 ),
( 4998 ),
( 5001 ),
( 5003 ),
( 5006 ),
( 5009 ),
( 5011 ),
( 5014 ),
( 5016 ),
( 5019 ),
( 5022 ),
( 5024 ),
( 5027 ),
( 5030 ),
( 5032 ),
( 5035 ),
( 5038 ),
( 5040 ),
( 5043 ),
( 5046 ),
( 5048 ),
( 5051 ),
( 5054 ),
( 5056 ),
( 5059 ),
( 5062 ),
( 5064 ),
( 5067 ),
( 5070 ),
( 5072 ),
( 5075 ),
( 5078 ),
( 5080 ),
( 5083 ),
( 5086 ),
( 5088 ),
( 5091 ),
( 5094 ),
( 5097 ),
( 5099 ),
( 5102 ),
( 5105 ),
( 5107 ),
( 5110 ),
( 5113 ),
( 5116 ),
( 5118 ),
( 5121 ),
( 5124 ),
( 5127 ),
( 5129 ),
( 5132 ),
( 5135 ),
( 5138 ),
( 5140 ),
( 5143 ),
( 5146 ),
( 5149 ),
( 5151 ),
( 5154 ),
( 5157 ),
( 5160 ),
( 5163 ),
( 5165 ),
( 5168 ),
( 5171 ),
( 5174 ),
( 5176 ),
( 5179 ),
( 5182 ),
( 5185 ),
( 5188 ),
( 5190 ),
( 5193 ),
( 5196 ),
( 5199 ),
( 5202 ),
( 5205 ),
( 5207 ),
( 5210 ),
( 5213 ),
( 5216 ),
( 5219 ),
( 5222 ),
( 5224 ),
( 5227 ),
( 5230 ),
( 5233 ),
( 5236 ),
( 5239 ),
( 5242 ),
( 5245 ),
( 5247 ),
( 5250 ),
( 5253 ),
( 5256 ),
( 5259 ),
( 5262 ),
( 5265 ),
( 5268 ),
( 5270 ),
( 5273 ),
( 5276 ),
( 5279 ),
( 5282 ),
( 5285 ),
( 5288 ),
( 5291 ),
( 5294 ),
( 5297 ),
( 5300 ),
( 5303 ),
( 5306 ),
( 5308 ),
( 5311 ),
( 5314 ),
( 5317 ),
( 5320 ),
( 5323 ),
( 5326 ),
( 5329 ),
( 5332 ),
( 5335 ),
( 5338 ),
( 5341 ),
( 5344 ),
( 5347 ),
( 5350 ),
( 5353 ),
( 5356 ),
( 5359 ),
( 5362 ),
( 5365 ),
( 5368 ),
( 5371 ),
( 5374 ),
( 5377 ),
( 5380 ),
( 5383 ),
( 5386 ),
( 5389 ),
( 5392 ),
( 5395 ),
( 5398 ),
( 5401 ),
( 5404 ),
( 5407 ),
( 5410 ),
( 5414 ),
( 5417 ),
( 5420 ),
( 5423 ),
( 5426 ),
( 5429 ),
( 5432 ),
( 5435 ),
( 5438 ),
( 5441 ),
( 5444 ),
( 5447 ),
( 5451 ),
( 5454 ),
( 5457 ),
( 5460 ),
( 5463 ),
( 5466 ),
( 5469 ),
( 5472 ),
( 5475 ),
( 5479 ),
( 5482 ),
( 5485 ),
( 5488 ),
( 5491 ),
( 5494 ),
( 5497 ),
( 5501 ),
( 5504 ),
( 5507 ),
( 5510 ),
( 5513 ),
( 5516 ),
( 5520 ),
( 5523 ),
( 5526 ),
( 5529 ),
( 5532 ),
( 5536 ),
( 5539 ),
( 5542 ),
( 5545 ),
( 5548 ),
( 5552 ),
( 5555 ),
( 5558 ),
( 5561 ),
( 5565 ),
( 5568 ),
( 5571 ),
( 5574 ),
( 5578 ),
( 5581 ),
( 5584 ),
( 5587 ),
( 5591 ),
( 5594 ),
( 5597 ),
( 5600 ),
( 5604 ),
( 5607 ),
( 5610 ),
( 5613 ),
( 5617 ),
( 5620 ),
( 5623 ),
( 5627 ),
( 5630 ),
( 5633 ),
( 5637 ),
( 5640 ),
( 5643 ),
( 5647 ),
( 5650 ),
( 5653 ),
( 5657 ),
( 5660 ),
( 5663 ),
( 5667 ),
( 5670 ),
( 5673 ),
( 5677 ),
( 5680 ),
( 5683 ),
( 5687 ),
( 5690 ),
( 5694 ),
( 5697 ),
( 5700 ),
( 5704 ),
( 5707 ),
( 5711 ),
( 5714 ),
( 5717 ),
( 5721 ),
( 5724 ),
( 5728 ),
( 5731 ),
( 5735 ),
( 5738 ),
( 5741 ),
( 5745 ),
( 5748 ),
( 5752 ),
( 5755 ),
( 5759 ),
( 5762 ),
( 5766 ),
( 5769 ),
( 5773 ),
( 5776 ),
( 5780 ),
( 5783 ),
( 5787 ),
( 5790 ),
( 5794 ),
( 5797 ),
( 5801 ),
( 5804 ),
( 5808 ),
( 5811 ),
( 5815 ),
( 5818 ),
( 5822 ),
( 5825 ),
( 5829 ),
( 5832 ),
( 5836 ),
( 5839 ),
( 5843 ),
( 5847 ),
( 5850 ),
( 5854 ),
( 5857 ),
( 5861 ),
( 5864 ),
( 5868 ),
( 5872 ),
( 5875 ),
( 5879 ),
( 5883 ),
( 5886 ),
( 5890 ),
( 5893 ),
( 5897 ),
( 5901 ),
( 5904 ),
( 5908 ),
( 5912 ),
( 5915 ),
( 5919 ),
( 5923 ),
( 5926 ),
( 5930 ),
( 5934 ),
( 5937 ),
( 5941 ),
( 5945 ),
( 5948 ),
( 5952 ),
( 5956 ),
( 5959 ),
( 5963 ),
( 5967 ),
( 5971 ),
( 5974 ),
( 5978 ),
( 5982 ),
( 5985 ),
( 5989 ),
( 5993 ),
( 5997 ),
( 6000 ),
( 6004 ),
( 6008 ),
( 6012 ),
( 6016 ),
( 6019 ),
( 6023 ),
( 6027 ),
( 6031 ),
( 6035 ),
( 6038 ),
( 6042 ),
( 6046 ),
( 6050 ),
( 6054 ),
( 6057 ),
( 6061 ),
( 6065 ),
( 6069 ),
( 6073 ),
( 6077 ),
( 6081 ),
( 6084 ),
( 6088 ),
( 6092 ),
( 6096 ),
( 6100 ),
( 6104 ),
( 6108 ),
( 6112 ),
( 6115 ),
( 6119 ),
( 6123 ),
( 6127 ),
( 6131 ),
( 6135 ),
( 6139 ),
( 6143 ),
( 6147 ),
( 6151 ),
( 6155 ),
( 6159 ),
( 6163 ),
( 6167 ),
( 6171 ),
( 6175 ),
( 6179 ),
( 6183 ),
( 6187 ),
( 6191 ),
( 6195 ),
( 6199 ),
( 6203 ),
( 6207 ),
( 6211 ),
( 6215 ),
( 6219 ),
( 6223 ),
( 6227 ),
( 6231 ),
( 6235 ),
( 6239 ),
( 6243 ),
( 6247 ),
( 6251 ),
( 6255 ),
( 6259 ),
( 6263 ),
( 6268 ),
( 6272 ),
( 6276 ),
( 6280 ),
( 6284 ),
( 6288 ),
( 6292 ),
( 6296 ),
( 6301 ),
( 6305 ),
( 6309 ),
( 6313 ),
( 6317 ),
( 6321 ),
( 6326 ),
( 6330 ),
( 6334 ),
( 6338 ),
( 6342 ),
( 6347 ),
( 6351 ),
( 6355 ),
( 6359 ),
( 6363 ),
( 6368 ),
( 6372 ),
( 6376 ),
( 6380 ),
( 6385 ),
( 6389 ),
( 6393 ),
( 6397 ),
( 6402 ),
( 6406 ),
( 6410 ),
( 6415 ),
( 6419 ),
( 6423 ),
( 6427 ),
( 6432 ),
( 6436 ),
( 6440 ),
( 6445 ),
( 6449 ),
( 6453 ),
( 6458 ),
( 6462 ),
( 6467 ),
( 6471 ),
( 6475 ),
( 6480 ),
( 6484 ),
( 6488 ),
( 6493 ),
( 6497 ),
( 6502 ),
( 6506 ),
( 6511 ),
( 6515 ),
( 6519 ),
( 6524 ),
( 6528 ),
( 6533 ),
( 6537 ),
( 6542 ),
( 6546 ),
( 6551 ),
( 6555 ),
( 6560 ),
( 6564 ),
( 6569 ),
( 6573 ),
( 6578 ),
( 6582 ),
( 6587 ),
( 6591 ),
( 6596 ),
( 6600 ),
( 6605 ),
( 6609 ),
( 6614 ),
( 6619 ),
( 6623 ),
( 6628 ),
( 6632 ),
( 6637 ),
( 6641 ),
( 6646 ),
( 6651 ),
( 6655 ),
( 6660 ),
( 6665 ),
( 6669 ),
( 6674 ),
( 6679 ),
( 6683 ),
( 6688 ),
( 6693 ),
( 6697 ),
( 6702 ),
( 6707 ),
( 6711 ),
( 6716 ),
( 6721 ),
( 6725 ),
( 6730 ),
( 6735 ),
( 6740 ),
( 6744 ),
( 6749 ),
( 6754 ),
( 6759 ),
( 6763 ),
( 6768 ),
( 6773 ),
( 6778 ),
( 6783 ),
( 6787 ),
( 6792 ),
( 6797 ),
( 6802 ),
( 6807 ),
( 6812 ),
( 6816 ),
( 6821 ),
( 6826 ),
( 6831 ),
( 6836 ),
( 6841 ),
( 6846 ),
( 6851 ),
( 6855 ),
( 6860 ),
( 6865 ),
( 6870 ),
( 6875 ),
( 6880 ),
( 6885 ),
( 6890 ),
( 6895 ),
( 6900 ),
( 6905 ),
( 6910 ),
( 6915 ),
( 6920 ),
( 6925 ),
( 6930 ),
( 6935 ),
( 6940 ),
( 6945 ),
( 6950 ),
( 6955 ),
( 6960 ),
( 6965 ),
( 6970 ),
( 6975 ),
( 6980 ),
( 6986 ),
( 6991 ),
( 6996 ),
( 7001 ),
( 7006 ),
( 7011 ),
( 7016 ),
( 7021 ),
( 7027 ),
( 7032 ),
( 7037 ),
( 7042 ),
( 7047 ),
( 7052 ),
( 7058 ),
( 7063 ),
( 7068 ),
( 7073 ),
( 7078 ),
( 7084 ),
( 7089 ),
( 7094 ),
( 7099 ),
( 7105 ),
( 7110 ),
( 7115 ),
( 7121 ),
( 7126 ),
( 7131 ),
( 7137 ),
( 7142 ),
( 7147 ),
( 7153 ),
( 7158 ),
( 7163 ),
( 7169 ),
( 7174 ),
( 7179 ),
( 7185 ),
( 7190 ),
( 7196 ),
( 7201 ),
( 7206 ),
( 7212 ),
( 7217 ),
( 7223 ),
( 7228 ),
( 7234 ),
( 7239 ),
( 7245 ),
( 7250 ),
( 7255 ),
( 7261 ),
( 7267 ),
( 7272 ),
( 7278 ),
( 7283 ),
( 7289 ),
( 7294 ),
( 7300 ),
( 7305 ),
( 7311 ),
( 7316 ),
( 7322 ),
( 7328 ),
( 7333 ),
( 7339 ),
( 7345 ),
( 7350 ),
( 7356 ),
( 7361 ),
( 7367 ),
( 7373 ),
( 7379 ),
( 7384 ),
( 7390 ),
( 7396 ),
( 7401 ),
( 7407 ),
( 7413 ),
( 7419 ),
( 7424 ),
( 7430 ),
( 7436 ),
( 7442 ),
( 7447 ),
( 7453 ),
( 7459 ),
( 7465 ),
( 7471 ),
( 7476 ),
( 7482 ),
( 7488 ),
( 7494 ),
( 7500 ),
( 7506 ),
( 7512 ),
( 7518 ),
( 7523 ),
( 7529 ),
( 7535 ),
( 7541 ),
( 7547 ),
( 7553 ),
( 7559 ),
( 7565 ),
( 7571 ),
( 7577 ),
( 7583 ),
( 7589 ),
( 7595 ),
( 7601 ),
( 7607 ),
( 7613 ),
( 7619 ),
( 7625 ),
( 7631 ),
( 7637 ),
( 7644 ),
( 7650 ),
( 7656 ),
( 7662 ),
( 7668 ),
( 7674 ),
( 7680 ),
( 7687 ),
( 7693 ),
( 7699 ),
( 7705 ),
( 7711 ),
( 7718 ),
( 7724 ),
( 7730 ),
( 7736 ),
( 7742 ),
( 7749 ),
( 7755 ),
( 7761 ),
( 7768 ),
( 7774 ),
( 7780 ),
( 7787 ),
( 7793 ),
( 7799 ),
( 7806 ),
( 7812 ),
( 7818 ),
( 7825 ),
( 7831 ),
( 7838 ),
( 7844 ),
( 7850 ),
( 7857 ),
( 7863 ),
( 7870 ),
( 7876 ),
( 7883 ),
( 7889 ),
( 7896 ),
( 7902 ),
( 7909 ),
( 7915 ),
( 7922 ),
( 7928 ),
( 7935 ),
( 7942 ),
( 7948 ),
( 7955 ),
( 7961 ),
( 7968 ),
( 7975 ),
( 7981 ),
( 7988 ),
( 7995 ),
( 8001 ),
( 8008 ),
( 8015 ),
( 8021 ),
( 8028 ),
( 8035 ),
( 8042 ),
( 8048 ),
( 8055 ),
( 8062 ),
( 8069 ),
( 8076 ),
( 8082 ),
( 8089 ),
( 8096 ),
( 8103 ),
( 8110 ),
( 8117 ),
( 8123 ),
( 8130 ),
( 8137 ),
( 8144 ),
( 8151 ),
( 8158 ),
( 8165 ),
( 8172 ),
( 8179 ),
( 8186 ),
( 8193 ),
( 8200 ),
( 8207 ),
( 8214 ),
( 8221 ),
( 8228 ),
( 8235 ),
( 8242 ),
( 8249 ),
( 8257 ),
( 8264 ),
( 8271 ),
( 8278 ),
( 8285 ),
( 8292 ),
( 8300 ),
( 8307 ),
( 8314 ),
( 8321 ),
( 8328 ),
( 8336 ),
( 8343 ),
( 8350 ),
( 8357 ),
( 8365 ),
( 8372 ),
( 8379 ),
( 8387 ),
( 8394 ),
( 8401 ),
( 8409 ),
( 8416 ),
( 8424 ),
( 8431 ),
( 8439 ),
( 8446 ),
( 8453 ),
( 8461 ),
( 8468 ),
( 8476 ),
( 8483 ),
( 8491 ),
( 8498 ),
( 8506 ),
( 8514 ),
( 8521 ),
( 8529 ),
( 8536 ),
( 8544 ),
( 8552 ),
( 8559 ),
( 8567 ),
( 8575 ),
( 8582 ),
( 8590 ),
( 8598 ),
( 8605 ),
( 8613 ),
( 8621 ),
( 8629 ),
( 8636 ),
( 8644 ),
( 8652 ),
( 8660 ),
( 8668 ),
( 8676 ),
( 8683 ),
( 8691 ),
( 8699 ),
( 8707 ),
( 8715 ),
( 8723 ),
( 8731 ),
( 8739 ),
( 8747 ),
( 8755 ),
( 8763 ),
( 8771 ),
( 8779 ),
( 8787 ),
( 8795 ),
( 8803 ),
( 8811 ),
( 8819 ),
( 8828 ),
( 8836 ),
( 8844 ),
( 8852 ),
( 8860 ),
( 8868 ),
( 8877 ),
( 8885 ),
( 8893 ),
( 8901 ),
( 8910 ),
( 8918 ),
( 8926 ),
( 8935 ),
( 8943 ),
( 8951 ),
( 8960 ),
( 8968 ),
( 8976 ),
( 8985 ),
( 8993 ),
( 9002 ),
( 9010 ),
( 9019 ),
( 9027 ),
( 9036 ),
( 9044 ),
( 9053 ),
( 9061 ),
( 9070 ),
( 9079 ),
( 9087 ),
( 9096 ),
( 9105 ),
( 9113 ),
( 9122 ),
( 9131 ),
( 9139 ),
( 9148 ),
( 9157 ),
( 9166 ),
( 9174 ),
( 9183 ),
( 9192 ),
( 9201 ),
( 9210 ),
( 9218 ),
( 9227 ),
( 9236 ),
( 9245 ),
( 9254 ),
( 9263 ),
( 9272 ),
( 9281 ),
( 9290 ),
( 9299 ),
( 9308 ),
( 9317 ),
( 9326 ),
( 9335 ),
( 9344 ),
( 9354 ),
( 9363 ),
( 9372 ),
( 9381 ),
( 9390 ),
( 9399 ),
( 9409 ),
( 9418 ),
( 9427 ),
( 9437 ),
( 9446 ),
( 9455 ),
( 9465 ),
( 9474 ),
( 9483 ),
( 9493 ),
( 9502 ),
( 9512 ),
( 9521 ),
( 9530 ),
( 9540 ),
( 9549 ),
( 9559 ),
( 9569 ),
( 9578 ),
( 9588 ),
( 9597 ),
( 9607 ),
( 9617 ),
( 9626 ),
( 9636 ),
( 9646 ),
( 9655 ),
( 9665 ),
( 9675 ),
( 9685 ),
( 9695 ),
( 9704 ),
( 9714 ),
( 9724 ),
( 9734 ),
( 9744 ),
( 9754 ),
( 9764 ),
( 9774 ),
( 9784 ),
( 9794 ),
( 9804 ),
( 9814 ),
( 9824 ),
( 9834 ),
( 9844 ),
( 9854 ),
( 9864 ),
( 9874 ),
( 9885 ),
( 9895 ),
( 9905 ),
( 9915 ),
( 9926 ),
( 9936 ),
( 9946 ),
( 9957 ),
( 9967 ),
( 9977 ),
( 9988 ),
( 9998 ),
( 10009 ),
( 10019 ),
( 10030 ),
( 10040 ),
( 10051 ),
( 10061 ),
( 10072 ),
( 10082 ),
( 10093 ),
( 10104 ),
( 10114 ),
( 10125 ),
( 10136 ),
( 10147 ),
( 10157 ),
( 10168 ),
( 10179 ),
( 10190 ),
( 10201 ),
( 10211 ),
( 10222 ),
( 10233 ),
( 10244 ),
( 10255 ),
( 10266 ),
( 10277 ),
( 10288 ),
( 10299 ),
( 10310 ),
( 10322 ),
( 10333 ),
( 10344 ),
( 10355 ),
( 10366 ),
( 10378 ),
( 10389 ),
( 10400 ),
( 10411 ),
( 10423 ),
( 10434 ),
( 10445 ),
( 10457 ),
( 10468 ),
( 10480 ),
( 10491 ),
( 10503 ),
( 10514 ),
( 10526 ),
( 10537 ),
( 10549 ),
( 10561 ),
( 10572 ),
( 10584 ),
( 10596 ),
( 10607 ),
( 10619 ),
( 10631 ),
( 10643 ),
( 10655 ),
( 10667 ),
( 10678 ),
( 10690 ),
( 10702 ),
( 10714 ),
( 10726 ),
( 10738 ),
( 10750 ),
( 10762 ),
( 10775 ),
( 10787 ),
( 10799 ),
( 10811 ),
( 10823 ),
( 10836 ),
( 10848 ),
( 10860 ),
( 10872 ),
( 10885 ),
( 10897 ),
( 10910 ),
( 10922 ),
( 10935 ),
( 10947 ),
( 10960 ),
( 10972 ),
( 10985 ),
( 10997 ),
( 11010 ),
( 11023 ),
( 11035 ),
( 11048 ),
( 11061 ),
( 11074 ),
( 11086 ),
( 11099 ),
( 11112 ),
( 11125 ),
( 11138 ),
( 11151 ),
( 11164 ),
( 11177 ),
( 11190 ),
( 11203 ),
( 11216 ),
( 11230 ),
( 11243 ),
( 11256 ),
( 11269 ),
( 11282 ),
( 11296 ),
( 11309 ),
( 11322 ),
( 11336 ),
( 11349 ),
( 11363 ),
( 11376 ),
( 11390 ),
( 11403 ),
( 11417 ),
( 11431 ),
( 11444 ),
( 11458 ),
( 11472 ),
( 11485 ),
( 11499 ),
( 11513 ),
( 11527 ),
( 11541 ),
( 11555 ),
( 11569 ),
( 11583 ),
( 11597 ),
( 11611 ),
( 11625 ),
( 11639 ),
( 11653 ),
( 11667 ),
( 11682 ),
( 11696 ),
( 11710 ),
( 11725 ),
( 11739 ),
( 11753 ),
( 11768 ),
( 11782 ),
( 11797 ),
( 11811 ),
( 11826 ),
( 11841 ),
( 11855 ),
( 11870 ),
( 11885 ),
( 11899 ),
( 11914 ),
( 11929 ),
( 11944 ),
( 11959 ),
( 11974 ),
( 11989 ),
( 12004 ),
( 12019 ),
( 12034 ),
( 12049 ),
( 12064 ),
( 12080 ),
( 12095 ),
( 12110 ),
( 12125 ),
( 12141 ),
( 12156 ),
( 12172 ),
( 12187 ),
( 12203 ),
( 12218 ),
( 12234 ),
( 12250 ),
( 12265 ),
( 12281 ),
( 12297 ),
( 12313 ),
( 12328 ),
( 12344 ),
( 12360 ),
( 12376 ),
( 12392 ),
( 12408 ),
( 12424 ),
( 12441 ),
( 12457 ),
( 12473 ),
( 12489 ),
( 12506 ),
( 12522 ),
( 12538 ),
( 12555 ),
( 12571 ),
( 12588 ),
( 12604 ),
( 12621 ),
( 12638 ),
( 12654 ),
( 12671 ),
( 12688 ),
( 12705 ),
( 12722 ),
( 12738 ),
( 12755 ),
( 12772 ),
( 12790 ),
( 12807 ),
( 12824 ),
( 12841 ),
( 12858 ),
( 12876 ),
( 12893 ),
( 12910 ),
( 12928 ),
( 12945 ),
( 12963 ),
( 12980 ),
( 12998 ),
( 13016 ),
( 13033 ),
( 13051 ),
( 13069 ),
( 13087 ),
( 13105 ),
( 13123 ),
( 13141 ),
( 13159 ),
( 13177 ),
( 13195 ),
( 13213 ),
( 13231 ),
( 13250 ),
( 13268 ),
( 13286 ),
( 13305 ),
( 13323 ),
( 13342 ),
( 13361 ),
( 13379 ),
( 13398 ),
( 13417 ),
( 13436 ),
( 13455 ),
( 13473 ),
( 13492 ),
( 13511 ),
( 13531 ),
( 13550 ),
( 13569 ),
( 13588 ),
( 13607 ),
( 13627 ),
( 13646 ),
( 13666 ),
( 13685 ),
( 13705 ),
( 13725 ),
( 13744 ),
( 13764 ),
( 13784 ),
( 13804 ),
( 13824 ),
( 13844 ),
( 13864 ),
( 13884 ),
( 13904 ),
( 13924 ),
( 13944 ),
( 13965 ),
( 13985 ),
( 14006 ),
( 14026 ),
( 14047 ),
( 14067 ),
( 14088 ),
( 14109 ),
( 14130 ),
( 14150 ),
( 14171 ),
( 14192 ),
( 14214 ),
( 14235 ),
( 14256 ),
( 14277 ),
( 14298 ),
( 14320 ),
( 14341 ),
( 14363 ),
( 14384 ),
( 14406 ),
( 14428 ),
( 14449 ),
( 14471 ),
( 14493 ),
( 14515 ),
( 14537 ),
( 14559 ),
( 14582 ),
( 14604 ),
( 14626 ),
( 14648 ),
( 14671 ),
( 14693 ),
( 14716 ),
( 14739 ),
( 14761 ),
( 14784 ),
( 14807 ),
( 14830 ),
( 14853 ),
( 14876 ),
( 14899 ),
( 14922 ),
( 14946 ),
( 14969 ),
( 14993 ),
( 15016 ),
( 15040 ),
( 15063 ),
( 15087 ),
( 15111 ),
( 15135 ),
( 15159 ),
( 15183 ),
( 15207 ),
( 15231 ),
( 15255 ),
( 15280 ),
( 15304 ),
( 15329 ),
( 15353 ),
( 15378 ),
( 15403 ),
( 15427 ),
( 15452 ),
( 15477 ),
( 15502 ),
( 15527 ),
( 15553 ),
( 15578 ),
( 15603 ),
( 15629 ),
( 15654 ),
( 15680 ),
( 15706 ),
( 15732 ),
( 15757 ),
( 15783 ),
( 15809 ),
( 15836 ),
( 15862 ),
( 15888 ),
( 15915 ),
( 15941 ),
( 15968 ),
( 15994 ),
( 16021 ),
( 16048 ),
( 16075 ),
( 16102 ),
( 16129 ),
( 16156 ),
( 16184 ),
( 16211 ),
( 16238 ),
( 16266 ),
( 16294 ),
( 16321 ),
( 16349 ),
( 16377 ),
( 16405 ),
( 16434 ),
( 16462 ),
( 16490 ),
( 16519 ),
( 16547 ),
( 16576 ),
( 16605 ),
( 16633 ),
( 16662 ),
( 16691 ),
( 16721 ),
( 16750 ),
( 16779 ),
( 16809 ),
( 16838 ),
( 16868 ),
( 16898 ),
( 16927 ),
( 16957 ),
( 16988 ),
( 17018 ),
( 17048 ),
( 17078 ),
( 17109 ),
( 17140 ),
( 17170 ),
( 17201 ),
( 17232 ),
( 17263 ),
( 17294 ),
( 17326 ),
( 17357 ),
( 17389 ),
( 17420 ),
( 17452 ),
( 17484 ),
( 17516 ),
( 17548 ),
( 17580 ),
( 17613 ),
( 17645 ),
( 17678 ),
( 17710 ),
( 17743 ),
( 17776 ),
( 17809 ),
( 17842 ),
( 17876 ),
( 17909 ),
( 17943 ),
( 17976 ),
( 18010 ),
( 18044 ),
( 18078 ),
( 18112 ),
( 18147 ),
( 18181 ),
( 18216 ),
( 18250 ),
( 18285 ),
( 18320 ),
( 18355 ),
( 18391 ),
( 18426 ),
( 18462 ),
( 18497 ),
( 18533 ),
( 18569 ),
( 18605 ),
( 18641 ),
( 18678 ),
( 18714 ),
( 18751 ),
( 18788 ),
( 18825 ),
( 18862 ),
( 18899 ),
( 18936 ),
( 18974 ),
( 19011 ),
( 19049 ),
( 19087 ),
( 19125 ),
( 19164 ),
( 19202 ),
( 19241 ),
( 19279 ),
( 19318 ),
( 19357 ),
( 19397 ),
( 19436 ),
( 19475 ),
( 19515 ),
( 19555 ),
( 19595 ),
( 19635 ),
( 19676 ),
( 19716 ),
( 19757 ),
( 19798 ),
( 19839 ),
( 19880 ),
( 19921 ),
( 19963 ),
( 20004 ),
( 20046 ),
( 20088 ),
( 20131 ),
( 20173 ),
( 20216 ),
( 20258 ),
( 20301 ),
( 20345 ),
( 20388 ),
( 20431 ),
( 20475 ),
( 20519 ),
( 20563 ),
( 20607 ),
( 20652 ),
( 20696 ),
( 20741 ),
( 20786 ),
( 20831 ),
( 20877 ),
( 20922 ),
( 20968 ),
( 21014 ),
( 21061 ),
( 21107 ),
( 21154 ),
( 21200 ),
( 21247 ),
( 21295 ),
( 21342 ),
( 21390 ),
( 21438 ),
( 21486 ),
( 21534 ),
( 21583 ),
( 21631 ),
( 21680 ),
( 21730 ),
( 21779 ),
( 21829 ),
( 21879 ),
( 21929 ),
( 21979 ),
( 22030 ),
( 22080 ),
( 22132 ),
( 22183 ),
( 22234 ),
( 22286 ),
( 22338 ),
( 22390 ),
( 22443 ),
( 22496 ),
( 22548 ),
( 22602 ),
( 22655 ),
( 22709 ),
( 22763 ),
( 22817 ),
( 22872 ),
( 22926 ),
( 22981 ),
( 23037 ),
( 23092 ),
( 23148 ),
( 23204 ),
( 23261 ),
( 23317 ),
( 23374 ),
( 23431 ),
( 23489 ),
( 23547 ),
( 23605 ),
( 23663 ),
( 23722 ),
( 23781 ),
( 23840 ),
( 23899 ),
( 23959 ),
( 24019 ),
( 24080 ),
( 24140 ),
( 24201 ),
( 24263 ),
( 24324 ),
( 24386 ),
( 24449 ),
( 24511 ),
( 24574 ),
( 24637 ),
( 24701 ),
( 24765 ),
( 24829 ),
( 24894 ),
( 24958 ),
( 25024 ),
( 25089 ),
( 25155 ),
( 25221 ),
( 25288 ),
( 25355 ),
( 25422 ),
( 25490 ),
( 25558 ),
( 25626 ),
( 25695 ),
( 25764 ),
( 25834 ),
( 25904 ),
( 25974 ),
( 26045 ),
( 26116 ),
( 26187 ),
( 26259 ),
( 26331 ),
( 26404 ),
( 26477 ),
( 26550 ),
( 26624 ),
( 26698 ),
( 26773 ),
( 26848 ),
( 26924 ),
( 26999 ),
( 27076 ),
( 27153 ),
( 27230 ),
( 27307 ),
( 27386 ),
( 27464 ),
( 27543 ),
( 27623 ),
( 27703 ),
( 27783 ),
( 27864 ),
( 27945 ),
( 28027 ),
( 28109 ),
( 28192 ),
( 28275 ),
( 28359 ),
( 28443 ),
( 28528 ),
( 28613 ),
( 28699 ),
( 28785 ),
( 28872 ),
( 28959 ),
( 29047 ),
( 29136 ),
( 29225 ),
( 29314 ),
( 29404 ),
( 29495 ),
( 29586 ),
( 29678 ),
( 29770 ),
( 29863 ),
( 29956 ),
( 30050 ),
( 30145 ),
( 30240 ),
( 30336 ),
( 30432 ),
( 30529 ),
( 30627 ),
( 30725 ),
( 30824 ),
( 30924 ),
( 31024 ),
( 31125 ),
( 31226 ),
( 31328 ),
( 31431 ),
( 31535 ),
( 31639 ),
( 31744 ),
( 31849 ),
( 31956 ),
( 32063 ),
( 32170 ),
( 32279 ),
( 32388 ),
( 32498 ),
( 32609 ),
( 32720 ),
( 32832 ),
( 32945 ),
( 33059 ),
( 33174 ),
( 33289 ),
( 33405 ),
( 33522 ),
( 33640 ),
( 33758 ),
( 33878 ),
( 33998 ),
( 34119 ),
( 34241 ),
( 34364 ),
( 34488 ),
( 34613 ),
( 34738 ),
( 34865 ),
( 34992 ),
( 35121 ),
( 35250 ),
( 35380 ),
( 35511 ),
( 35644 ),
( 35777 ),
( 35911 ),
( 36046 ),
( 36182 ),
( 36320 ),
( 36458 ),
( 36597 ),
( 36738 ),
( 36879 ),
( 37022 ),
( 37166 ),
( 37310 ),
( 37456 ),
( 37603 ),
( 37752 ),
( 37901 ),
( 38052 ),
( 38204 ),
( 38357 ),
( 38511 ),
( 38666 ),
( 38823 ),
( 38981 ),
( 39141 ),
( 39301 ),
( 39463 ),
( 39627 ),
( 39791 ),
( 39957 ),
( 40125 ),
( 40294 ),
( 40464 ),
( 40636 ),
( 40809 ),
( 40984 ),
( 41160 ),
( 41337 ),
( 41517 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 ),
( 41666 )
);




end package LUT_pkg;
