library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (
(	7049	)	,
(	7034	)	,
(	7019	)	,
(	7004	)	,
(	6989	)	,
(	6974	)	,
(	6959	)	,
(	6944	)	,
(	6929	)	,
(	6914	)	,
(	6900	)	,
(	6885	)	,
(	6870	)	,
(	6855	)	,
(	6841	)	,
(	6826	)	,
(	6811	)	,
(	6797	)	,
(	6782	)	,
(	6767	)	,
(	6753	)	,
(	6738	)	,
(	6724	)	,
(	6710	)	,
(	6695	)	,
(	6681	)	,
(	6666	)	,
(	6652	)	,
(	6638	)	,
(	6623	)	,
(	6609	)	,
(	6595	)	,
(	6581	)	,
(	6567	)	,
(	6552	)	,
(	6538	)	,
(	6524	)	,
(	6510	)	,
(	6496	)	,
(	6482	)	,
(	6468	)	,
(	6454	)	,
(	6440	)	,
(	6426	)	,
(	6413	)	,
(	6399	)	,
(	6385	)	,
(	6371	)	,
(	6357	)	,
(	6344	)	,
(	6330	)	,
(	6316	)	,
(	6303	)	,
(	6289	)	,
(	6275	)	,
(	6262	)	,
(	6248	)	,
(	6235	)	,
(	6221	)	,
(	6208	)	,
(	6194	)	,
(	6181	)	,
(	6167	)	,
(	6154	)	,
(	6141	)	,
(	6127	)	,
(	6114	)	,
(	6101	)	,
(	6088	)	,
(	6074	)	,
(	6061	)	,
(	6048	)	,
(	6035	)	,
(	6022	)	,
(	6009	)	,
(	5996	)	,
(	5983	)	,
(	5970	)	,
(	5957	)	,
(	5944	)	,
(	5931	)	,
(	5918	)	,
(	5905	)	,
(	5892	)	,
(	5879	)	,
(	5867	)	,
(	5854	)	,
(	5841	)	,
(	5828	)	,
(	5816	)	,
(	5803	)	,
(	5790	)	,
(	5778	)	,
(	5765	)	,
(	5753	)	,
(	5740	)	,
(	5728	)	,
(	5715	)	,
(	5703	)	,
(	5690	)	,
(	5678	)	,
(	5665	)	,
(	5653	)	,
(	5641	)	,
(	5628	)	,
(	5616	)	,
(	5604	)	,
(	5592	)	,
(	5579	)	,
(	5567	)	,
(	5555	)	,
(	5543	)	,
(	5531	)	,
(	5519	)	,
(	5507	)	,
(	5495	)	,
(	5483	)	,
(	5471	)	,
(	5459	)	,
(	5447	)	,
(	5435	)	,
(	5423	)	,
(	5411	)	,
(	5399	)	,
(	5387	)	,
(	5376	)	,
(	5364	)	,
(	5352	)	,
(	5340	)	,
(	5329	)	,
(	5317	)	,
(	5305	)	,
(	5294	)	,
(	5282	)	,
(	5270	)	,
(	5259	)	,
(	5247	)	,
(	5236	)	,
(	5224	)	,
(	5213	)	,
(	5201	)	,
(	5190	)	,
(	5179	)	,
(	5167	)	,
(	5156	)	,
(	5145	)	,
(	5133	)	,
(	5122	)	,
(	5111	)	,
(	5100	)	,
(	5088	)	,
(	5077	)	,
(	5066	)	,
(	5055	)	,
(	5044	)	,
(	5033	)	,
(	5022	)	,
(	5011	)	,
(	5000	)	,
(	4989	)	,
(	4978	)	,
(	4967	)	,
(	4956	)	,
(	4945	)	,
(	4934	)	,
(	4923	)	,
(	4912	)	,
(	4902	)	,
(	4891	)	,
(	4880	)	,
(	4869	)	,
(	4859	)	,
(	4848	)	,
(	4837	)	,
(	4827	)	,
(	4816	)	,
(	4805	)	,
(	4795	)	,
(	4784	)	,
(	4774	)	,
(	4763	)	,
(	4753	)	,
(	4742	)	,
(	4732	)	,
(	4721	)	,
(	4711	)	,
(	4700	)	,
(	4690	)	,
(	4680	)	,
(	4669	)	,
(	4659	)	,
(	4649	)	,
(	4639	)	,
(	4628	)	,
(	4618	)	,
(	4608	)	,
(	4598	)	,
(	4588	)	,
(	4578	)	,
(	4568	)	,
(	4557	)	,
(	4547	)	,
(	4537	)	,
(	4527	)	,
(	4517	)	,
(	4507	)	,
(	4498	)	,
(	4488	)	,
(	4478	)	,
(	4468	)	,
(	4458	)	,
(	4448	)	,
(	4438	)	,
(	4429	)	,
(	4419	)	,
(	4409	)	,
(	4399	)	,
(	4390	)	,
(	4380	)	,
(	4370	)	,
(	4361	)	,
(	4351	)	,
(	4341	)	,
(	4332	)	,
(	4322	)	,
(	4313	)	,
(	4303	)	,
(	4294	)	,
(	4284	)	,
(	4275	)	,
(	4265	)	,
(	4256	)	,
(	4246	)	,
(	4237	)	,
(	4228	)	,
(	4218	)	,
(	4209	)	,
(	4200	)	,
(	4191	)	,
(	4181	)	,
(	4172	)	,
(	4163	)	,
(	4154	)	,
(	4145	)	,
(	4135	)	,
(	4126	)	,
(	4117	)	,
(	4108	)	,
(	4099	)	,
(	4090	)	,
(	4081	)	,
(	4072	)	,
(	4063	)	,
(	4054	)	,
(	4045	)	,
(	4036	)	,
(	4027	)	,
(	4018	)	,
(	4009	)	,
(	4001	)	,
(	3992	)	,
(	3983	)	,
(	3974	)	,
(	3965	)	,
(	3957	)	,
(	3948	)	,
(	3939	)	,
(	3931	)	,
(	3922	)	,
(	3913	)	,
(	3905	)	,
(	3896	)	,
(	3887	)	,
(	3879	)	,
(	3870	)	,
(	3862	)	,
(	3853	)	,
(	3845	)	,
(	3836	)	,
(	3828	)	,
(	3819	)	,
(	3811	)	,
(	3803	)	,
(	3794	)	,
(	3786	)	,
(	3778	)	,
(	3769	)	,
(	3761	)	,
(	3753	)	,
(	3744	)	,
(	3736	)	,
(	3728	)	,
(	3720	)	,
(	3712	)	,
(	3703	)	,
(	3695	)	,
(	3687	)	,
(	3679	)	,
(	3671	)	,
(	3663	)	,
(	3655	)	,
(	3647	)	,
(	3639	)	,
(	3631	)	,
(	3623	)	,
(	3615	)	,
(	3607	)	,
(	3599	)	,
(	3591	)	,
(	3583	)	,
(	3575	)	,
(	3567	)	,
(	3560	)	,
(	3552	)	,
(	3544	)	,
(	3536	)	,
(	3528	)	,
(	3521	)	,
(	3513	)	,
(	3505	)	,
(	3498	)	,
(	3490	)	,
(	3482	)	,
(	3475	)	,
(	3467	)	,
(	3459	)	,
(	3452	)	,
(	3444	)	,
(	3437	)	,
(	3429	)	,
(	3422	)	,
(	3414	)	,
(	3407	)	,
(	3399	)	,
(	3392	)	,
(	3384	)	,
(	3377	)	,
(	3370	)	,
(	3362	)	,
(	3355	)	,
(	3348	)	,
(	3340	)	,
(	3333	)	,
(	3326	)	,
(	3319	)	,
(	3311	)	,
(	3304	)	,
(	3297	)	,
(	3290	)	,
(	3282	)	,
(	3275	)	,
(	3268	)	,
(	3261	)	,
(	3254	)	,
(	3247	)	,
(	3240	)	,
(	3233	)	,
(	3226	)	,
(	3219	)	,
(	3212	)	,
(	3205	)	,
(	3198	)	,
(	3191	)	,
(	3184	)	,
(	3177	)	,
(	3170	)	,
(	3163	)	,
(	3156	)	,
(	3149	)	,
(	3143	)	,
(	3136	)	,
(	3129	)	,
(	3122	)	,
(	3115	)	,
(	3109	)	,
(	3102	)	,
(	3095	)	,
(	3089	)	,
(	3082	)	,
(	3075	)	,
(	3069	)	,
(	3062	)	,
(	3055	)	,
(	3049	)	,
(	3042	)	,
(	3035	)	,
(	3029	)	,
(	3022	)	,
(	3016	)	,
(	3009	)	,
(	3003	)	,
(	2996	)	,
(	2990	)	,
(	2984	)	,
(	2977	)	,
(	2971	)	,
(	2964	)	,
(	2958	)	,
(	2952	)	,
(	2945	)	,
(	2939	)	,
(	2933	)	,
(	2926	)	,
(	2920	)	,
(	2914	)	,
(	2907	)	,
(	2901	)	,
(	2895	)	,
(	2889	)	,
(	2883	)	,
(	2876	)	,
(	2870	)	,
(	2864	)	,
(	2858	)	,
(	2852	)	,
(	2846	)	,
(	2840	)	,
(	2834	)	,
(	2828	)	,
(	2822	)	,
(	2816	)	,
(	2810	)	,
(	2804	)	,
(	2798	)	,
(	2792	)	,
(	2786	)	,
(	2780	)	,
(	2774	)	,
(	2768	)	,
(	2762	)	,
(	2756	)	,
(	2750	)	,
(	2744	)	,
(	2739	)	,
(	2733	)	,
(	2727	)	,
(	2721	)	,
(	2715	)	,
(	2710	)	,
(	2704	)	,
(	2698	)	,
(	2693	)	,
(	2687	)	,
(	2681	)	,
(	2676	)	,
(	2670	)	,
(	2664	)	,
(	2659	)	,
(	2653	)	,
(	2647	)	,
(	2642	)	,
(	2636	)	,
(	2631	)	,
(	2625	)	,
(	2620	)	,
(	2614	)	,
(	2609	)	,
(	2603	)	,
(	2598	)	,
(	2592	)	,
(	2587	)	,
(	2581	)	,
(	2576	)	,
(	2571	)	,
(	2565	)	,
(	2560	)	,
(	2555	)	,
(	2549	)	,
(	2544	)	,
(	2539	)	,
(	2533	)	,
(	2528	)	,
(	2523	)	,
(	2518	)	,
(	2512	)	,
(	2507	)	,
(	2502	)	,
(	2497	)	,
(	2492	)	,
(	2486	)	,
(	2481	)	,
(	2476	)	,
(	2471	)	,
(	2466	)	,
(	2461	)	,
(	2456	)	,
(	2451	)	,
(	2446	)	,
(	2440	)	,
(	2435	)	,
(	2430	)	,
(	2425	)	,
(	2420	)	,
(	2415	)	,
(	2411	)	,
(	2406	)	,
(	2401	)	,
(	2396	)	,
(	2391	)	,
(	2386	)	,
(	2381	)	,
(	2376	)	,
(	2371	)	,
(	2366	)	,
(	2362	)	,
(	2357	)	,
(	2352	)	,
(	2347	)	,
(	2342	)	,
(	2338	)	,
(	2333	)	,
(	2328	)	,
(	2323	)	,
(	2319	)	,
(	2314	)	,
(	2309	)	,
(	2305	)	,
(	2300	)	,
(	2295	)	,
(	2291	)	,
(	2286	)	,
(	2281	)	,
(	2277	)	,
(	2272	)	,
(	2268	)	,
(	2263	)	,
(	2259	)	,
(	2254	)	,
(	2249	)	,
(	2245	)	,
(	2240	)	,
(	2236	)	,
(	2232	)	,
(	2227	)	,
(	2223	)	,
(	2218	)	,
(	2214	)	,
(	2209	)	,
(	2205	)	,
(	2201	)	,
(	2196	)	,
(	2192	)	,
(	2187	)	,
(	2183	)	,
(	2179	)	,
(	2174	)	,
(	2170	)	,
(	2166	)	,
(	2162	)	,
(	2157	)	,
(	2153	)	,
(	2149	)	,
(	2145	)	,
(	2140	)	,
(	2136	)	,
(	2132	)	,
(	2128	)	,
(	2124	)	,
(	2119	)	,
(	2115	)	,
(	2111	)	,
(	2107	)	,
(	2103	)	,
(	2099	)	,
(	2095	)	,
(	2091	)	,
(	2087	)	,
(	2082	)	,
(	2078	)	,
(	2074	)	,
(	2070	)	,
(	2066	)	,
(	2062	)	,
(	2058	)	,
(	2054	)	,
(	2050	)	,
(	2046	)	,
(	2043	)	,
(	2039	)	,
(	2035	)	,
(	2031	)	,
(	2027	)	,
(	2023	)	,
(	2019	)	,
(	2015	)	,
(	2011	)	,
(	2008	)	,
(	2004	)	,
(	2000	)	,
(	1996	)	,
(	1992	)	,
(	1988	)	,
(	1985	)	,
(	1981	)	,
(	1977	)	,
(	1973	)	,
(	1970	)	,
(	1966	)	,
(	1962	)	,
(	1959	)	,
(	1955	)	,
(	1951	)	,
(	1948	)	,
(	1944	)	,
(	1940	)	,
(	1937	)	,
(	1933	)	,
(	1929	)	,
(	1926	)	,
(	1922	)	,
(	1919	)	,
(	1915	)	,
(	1911	)	,
(	1908	)	,
(	1904	)	,
(	1901	)	,
(	1897	)	,
(	1894	)	,
(	1890	)	,
(	1887	)	,
(	1883	)	,
(	1880	)	,
(	1876	)	,
(	1873	)	,
(	1869	)	,
(	1866	)	,
(	1863	)	,
(	1859	)	,
(	1856	)	,
(	1852	)	,
(	1849	)	,
(	1846	)	,
(	1842	)	,
(	1839	)	,
(	1836	)	,
(	1832	)	,
(	1829	)	,
(	1826	)	,
(	1822	)	,
(	1819	)	,
(	1816	)	,
(	1813	)	,
(	1809	)	,
(	1806	)	,
(	1803	)	,
(	1800	)	,
(	1796	)	,
(	1793	)	,
(	1790	)	,
(	1787	)	,
(	1784	)	,
(	1780	)	,
(	1777	)	,
(	1774	)	,
(	1771	)	,
(	1768	)	,
(	1765	)	,
(	1762	)	,
(	1758	)	,
(	1755	)	,
(	1752	)	,
(	1749	)	,
(	1746	)	,
(	1743	)	,
(	1740	)	,
(	1737	)	,
(	1734	)	,
(	1731	)	,
(	1728	)	,
(	1725	)	,
(	1722	)	,
(	1719	)	,
(	1716	)	,
(	1713	)	,
(	1710	)	,
(	1707	)	,
(	1704	)	,
(	1701	)	,
(	1698	)	,
(	1695	)	,
(	1693	)	,
(	1690	)	,
(	1687	)	,
(	1684	)	,
(	1681	)	,
(	1678	)	,
(	1675	)	,
(	1672	)	,
(	1670	)	,
(	1667	)	,
(	1664	)	,
(	1661	)	,
(	1658	)	,
(	1656	)	,
(	1653	)	,
(	1650	)	,
(	1647	)	,
(	1645	)	,
(	1642	)	,
(	1639	)	,
(	1636	)	,
(	1634	)	,
(	1631	)	,
(	1628	)	,
(	1626	)	,
(	1623	)	,
(	1620	)	,
(	1617	)	,
(	1615	)	,
(	1612	)	,
(	1610	)	,
(	1607	)	,
(	1604	)	,
(	1602	)	,
(	1599	)	,
(	1596	)	,
(	1594	)	,
(	1591	)	,
(	1589	)	,
(	1586	)	,
(	1584	)	,
(	1581	)	,
(	1578	)	,
(	1576	)	,
(	1573	)	,
(	1571	)	,
(	1568	)	,
(	1566	)	,
(	1563	)	,
(	1561	)	,
(	1558	)	,
(	1556	)	,
(	1553	)	,
(	1551	)	,
(	1549	)	,
(	1546	)	,
(	1544	)	,
(	1541	)	,
(	1539	)	,
(	1536	)	,
(	1534	)	,
(	1532	)	,
(	1529	)	,
(	1527	)	,
(	1525	)	,
(	1522	)	,
(	1520	)	,
(	1517	)	,
(	1515	)	,
(	1513	)	,
(	1510	)	,
(	1508	)	,
(	1506	)	,
(	1504	)	,
(	1501	)	,
(	1499	)	,
(	1497	)	,
(	1494	)	,
(	1492	)	,
(	1490	)	,
(	1488	)	,
(	1485	)	,
(	1483	)	,
(	1481	)	,
(	1479	)	,
(	1477	)	,
(	1474	)	,
(	1472	)	,
(	1470	)	,
(	1468	)	,
(	1466	)	,
(	1463	)	,
(	1461	)	,
(	1459	)	,
(	1457	)	,
(	1455	)	,
(	1453	)	,
(	1451	)	,
(	1448	)	,
(	1446	)	,
(	1444	)	,
(	1442	)	,
(	1440	)	,
(	1438	)	,
(	1436	)	,
(	1434	)	,
(	1432	)	,
(	1430	)	,
(	1428	)	,
(	1426	)	,
(	1424	)	,
(	1421	)	,
(	1419	)	,
(	1417	)	,
(	1415	)	,
(	1413	)	,
(	1411	)	,
(	1409	)	,
(	1407	)	,
(	1405	)	,
(	1404	)	,
(	1402	)	,
(	1400	)	,
(	1398	)	,
(	1396	)	,
(	1394	)	,
(	1392	)	,
(	1390	)	,
(	1388	)	,
(	1386	)	,
(	1384	)	,
(	1382	)	,
(	1380	)	,
(	1378	)	,
(	1377	)	,
(	1375	)	,
(	1373	)	,
(	1371	)	,
(	1369	)	,
(	1367	)	,
(	1365	)	,
(	1364	)	,
(	1362	)	,
(	1360	)	,
(	1358	)	,
(	1356	)	,
(	1355	)	,
(	1353	)	,
(	1351	)	,
(	1349	)	,
(	1347	)	,
(	1346	)	,
(	1344	)	,
(	1342	)	,
(	1340	)	,
(	1339	)	,
(	1337	)	,
(	1335	)	,
(	1333	)	,
(	1332	)	,
(	1330	)	,
(	1328	)	,
(	1326	)	,
(	1325	)	,
(	1323	)	,
(	1321	)	,
(	1320	)	,
(	1318	)	,
(	1316	)	,
(	1315	)	,
(	1313	)	,
(	1311	)	,
(	1310	)	,
(	1308	)	,
(	1306	)	,
(	1305	)	,
(	1303	)	,
(	1302	)	,
(	1300	)	,
(	1298	)	,
(	1297	)	,
(	1295	)	,
(	1294	)	,
(	1292	)	,
(	1290	)	,
(	1289	)	,
(	1287	)	,
(	1286	)	,
(	1284	)	,
(	1283	)	,
(	1281	)	,
(	1279	)	,
(	1278	)	,
(	1276	)	,
(	1275	)	,
(	1273	)	,
(	1272	)	,
(	1270	)	,
(	1269	)	,
(	1267	)	,
(	1266	)	,
(	1264	)	,
(	1263	)	,
(	1261	)	,
(	1260	)	,
(	1258	)	,
(	1257	)	,
(	1255	)	,
(	1254	)	,
(	1252	)	,
(	1251	)	,
(	1250	)	,
(	1248	)	,
(	1247	)	,
(	1245	)	,
(	1244	)	,
(	1242	)	,
(	1241	)	,
(	1240	)	,
(	1238	)	,
(	1237	)	,
(	1235	)	,
(	1234	)	,
(	1233	)	,
(	1231	)	,
(	1230	)	,
(	1229	)	,
(	1227	)	,
(	1226	)	,
(	1224	)	,
(	1223	)	,
(	1222	)	,
(	1220	)	,
(	1219	)	,
(	1218	)	,
(	1216	)	,
(	1215	)	,
(	1214	)	,
(	1212	)	,
(	1211	)	,
(	1210	)	,
(	1209	)	,
(	1207	)	,
(	1206	)	,
(	1205	)	,
(	1203	)	,
(	1202	)	,
(	1201	)	,
(	1200	)	,
(	1198	)	,
(	1197	)	,
(	1196	)	,
(	1195	)	,
(	1193	)	,
(	1192	)	,
(	1191	)	,
(	1190	)	,
(	1188	)	,
(	1187	)	,
(	1186	)	,
(	1185	)	,
(	1183	)	,
(	1182	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1177	)	,
(	1176	)	,
(	1175	)	,
(	1174	)	,
(	1173	)	,
(	1172	)	,
(	1170	)	,
(	1169	)	,
(	1168	)	,
(	1167	)	,
(	1166	)	,
(	1165	)	,
(	1163	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1159	)	,
(	1158	)	,
(	1157	)	,
(	1156	)	,
(	1154	)	,
(	1153	)	,
(	1152	)	,
(	1151	)	,
(	1150	)	,
(	1149	)	,
(	1148	)	,
(	1147	)	,
(	1146	)	,
(	1145	)	,
(	1144	)	,
(	1142	)	,
(	1141	)	,
(	1140	)	,
(	1139	)	,
(	1138	)	,
(	1137	)	,
(	1136	)	,
(	1135	)	,
(	1134	)	,
(	1133	)	,
(	1132	)	,
(	1131	)	,
(	1130	)	,
(	1129	)	,
(	1128	)	,
(	1127	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1121	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1116	)	,
(	1115	)	,
(	1114	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1105	)	,
(	1104	)	,
(	1103	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1099	)	,
(	1098	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1092	)	,
(	1091	)	,
(	1090	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1080	)	,
(	1079	)	,
(	1078	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1073	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1068	)	,
(	1068	)	,
(	1067	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1052	)	,
(	1052	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1032	)	,
(	1031	)	,
(	1030	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1027	)	,
(	1026	)	,
(	1025	)	,
(	1025	)	,
(	1024	)	,
(	1023	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1021	)	,
(	1020	)	,
(	1019	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1007	)	,
(	1006	)	,
(	1005	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1003	)	,
(	1002	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	1000	)	,
(	999	)	,
(	998	)	,
(	998	)	,
(	997	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	993	)	,
(	992	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	990	)	,
(	989	)	,
(	989	)	,
(	988	)	,
(	987	)	,
(	987	)	,
(	986	)	,
(	986	)	,
(	985	)	,
(	984	)	,
(	984	)	,
(	983	)	,
(	983	)	,
(	982	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	980	)	,
(	979	)	,
(	979	)	,
(	978	)	,
(	977	)	,
(	977	)	,
(	976	)	,
(	976	)	,
(	975	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	973	)	,
(	972	)	,
(	972	)	,
(	971	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	969	)	,
(	968	)	,
(	968	)	,
(	967	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	965	)	,
(	964	)	,
(	964	)	,
(	963	)	,
(	963	)	,
(	962	)	,
(	962	)	,
(	961	)	,
(	960	)	,
(	960	)	,
(	959	)	,
(	959	)	,
(	958	)	,
(	958	)	,
(	957	)	,
(	957	)	,
(	956	)	,
(	956	)	,
(	955	)	,
(	954	)	,
(	954	)	,
(	953	)	,
(	953	)	,
(	952	)	,
(	952	)	,
(	951	)	,
(	951	)	,
(	950	)	,
(	950	)	,
(	949	)	,
(	949	)	,
(	948	)	,
(	948	)	,
(	947	)	,
(	946	)	,
(	946	)	,
(	945	)	,
(	945	)	,
(	944	)	,
(	944	)	,
(	943	)	,
(	943	)	,
(	942	)	,
(	942	)	,
(	941	)	,
(	941	)	,
(	940	)	,
(	940	)	,
(	939	)	,
(	939	)	,
(	938	)	,
(	937	)	,
(	937	)	,
(	936	)	,
(	936	)	,
(	935	)	,
(	935	)	,
(	934	)	,
(	934	)	,
(	933	)	,
(	933	)	,
(	932	)	,
(	932	)	,
(	931	)	,
(	931	)	,
(	930	)	,
(	930	)	,
(	929	)	,
(	929	)	,
(	928	)	,
(	928	)	,
(	927	)	,
(	927	)	,
(	926	)	,
(	926	)	,
(	925	)	,
(	925	)	,
(	924	)	,
(	924	)	,
(	923	)	,
(	922	)	,
(	922	)	,
(	921	)	,
(	921	)	,
(	920	)	,
(	920	)	,
(	919	)	,
(	919	)	,
(	918	)	,
(	918	)	,
(	917	)	,
(	917	)	,
(	916	)	,
(	916	)	,
(	915	)	,
(	915	)	,
(	914	)	,
(	914	)	,
(	913	)	,
(	913	)	,
(	912	)	,
(	912	)	,
(	911	)	,
(	911	)	,
(	910	)	,
(	910	)	,
(	909	)	,
(	909	)	,
(	908	)	,
(	908	)	,
(	907	)	,
(	907	)	,
(	906	)	,
(	906	)	,
(	905	)	,
(	905	)	,
(	904	)	,
(	904	)	,
(	903	)	,
(	903	)	,
(	902	)	,
(	902	)	,
(	901	)	,
(	901	)	,
(	900	)	,
(	900	)	,
(	899	)	,
(	899	)	,
(	898	)	,
(	898	)	,
(	897	)	,
(	896	)	,
(	896	)	,
(	895	)	,
(	895	)	,
(	894	)	,
(	894	)	,
(	893	)	,
(	893	)	,
(	892	)	,
(	892	)	,
(	891	)	,
(	891	)	,
(	890	)	,
(	890	)	,
(	889	)	,
(	889	)	,
(	888	)	,
(	888	)	,
(	887	)	,
(	887	)	,
(	886	)	,
(	886	)	,
(	885	)	,
(	885	)	,
(	884	)	,
(	884	)	,
(	883	)	,
(	883	)	,
(	882	)	,
(	882	)	,
(	881	)	,
(	881	)	,
(	880	)	,
(	880	)	,
(	879	)	,
(	879	)	,
(	878	)	,
(	878	)	,
(	877	)	,
(	876	)	,
(	876	)	,
(	875	)	,
(	875	)	,
(	874	)	,
(	874	)	,
(	873	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	869	)	,
(	868	)	,
(	868	)	,
(	867	)	,
(	867	)	,
(	866	)	,
(	866	)	,
(	865	)	,
(	864	)	,
(	864	)	,
(	863	)	,
(	863	)	,
(	862	)	,
(	862	)	,
(	861	)	,
(	861	)	,
(	860	)	,
(	860	)	,
(	859	)	,
(	859	)	,
(	858	)	,
(	858	)	,
(	857	)	,
(	856	)	,
(	856	)	,
(	855	)	,
(	855	)	,
(	854	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	852	)	,
(	851	)	,
(	851	)	,
(	850	)	,
(	849	)	,
(	849	)	,
(	848	)	,
(	848	)	,
(	847	)	,
(	847	)	,
(	846	)	,
(	846	)	,
(	845	)	,
(	845	)	,
(	844	)	,
(	843	)	,
(	843	)	,
(	842	)	,
(	842	)	,
(	841	)	,
(	841	)	,
(	840	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	837	)	,
(	837	)	,
(	836	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	834	)	,
(	833	)	,
(	832	)	,
(	832	)	,
(	831	)	,
(	831	)	,
(	830	)	,
(	830	)	,
(	829	)	,
(	828	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	826	)	,
(	825	)	,
(	824	)	,
(	824	)	,
(	823	)	,
(	823	)	,
(	822	)	,
(	822	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	816	)	,
(	816	)	,
(	815	)	,
(	815	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	812	)	,
(	811	)	,
(	810	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	808	)	,
(	807	)	,
(	806	)	,
(	806	)	,
(	805	)	,
(	805	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	802	)	,
(	801	)	,
(	800	)	,
(	800	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	797	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	794	)	,
(	793	)	,
(	792	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	789	)	,
(	789	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	782	)	,
(	782	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	779	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	775	)	,
(	775	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	754	)	,
(	754	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	748	)	,
(	748	)	,
(	747	)	,
(	746	)	,
(	746	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	742	)	,
(	741	)	,
(	741	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	730	)	,
(	730	)	,
(	729	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	723	)	,
(	722	)	,
(	722	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	696	)	,
(	695	)	,
(	695	)	,
(	694	)	,
(	693	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	680	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	673	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	666	)	,
(	665	)	,
(	664	)	,
(	664	)	,
(	663	)	,
(	662	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	655	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	651	)	,
(	650	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	646	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	642	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	638	)	,
(	637	)	,
(	636	)	,
(	635	)	,
(	635	)	,
(	634	)	,
(	633	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	629	)	,
(	628	)	,
(	627	)	,
(	626	)	,
(	626	)	,
(	625	)	,
(	624	)	,
(	623	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	619	)	,
(	618	)	,
(	617	)	,
(	616	)	,
(	616	)	,
(	615	)	,
(	614	)	,
(	613	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	609	)	,
(	608	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	604	)	,
(	603	)	,
(	602	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	598	)	,
(	597	)	,
(	596	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	592	)	,
(	591	)	,
(	590	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	586	)	,
(	585	)	,
(	584	)	,
(	583	)	,
(	582	)	,
(	582	)	,
(	581	)	,
(	580	)	,
(	579	)	,
(	578	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	574	)	,
(	573	)	,
(	572	)	,
(	571	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	567	)	,
(	566	)	,
(	565	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	561	)	,
(	560	)	,
(	559	)	,
(	558	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	554	)	,
(	553	)	,
(	552	)	,
(	551	)	,
(	550	)	,
(	549	)	,
(	548	)	,
(	548	)	,
(	547	)	,
(	546	)	,
(	545	)	,
(	544	)	,
(	543	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	539	)	,
(	538	)	,
(	537	)	,
(	536	)	,
(	535	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	531	)	,
(	530	)	,
(	529	)	,
(	528	)	,
(	527	)	,
(	526	)	,
(	526	)	,
(	525	)	,
(	524	)	,
(	523	)	,
(	522	)	,
(	521	)	,
(	520	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	516	)	,
(	515	)	,
(	514	)	,
(	513	)	,
(	512	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	508	)	,
(	507	)	,
(	506	)	,
(	505	)	,
(	504	)	,
(	503	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	499	)	,
(	498	)	,
(	497	)	,
(	496	)	,
(	495	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	491	)	,
(	490	)	,
(	489	)	,
(	488	)	,
(	487	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	483	)	,
(	482	)	,
(	481	)	,
(	480	)	,
(	479	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	475	)	,
(	474	)	,
(	473	)	,
(	472	)	,
(	471	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	467	)	,
(	466	)	,
(	465	)	,
(	464	)	,
(	463	)	,
(	462	)	,
(	461	)	,
(	461	)	,
(	460	)	,
(	459	)	,
(	458	)	,
(	457	)	,
(	456	)	,
(	455	)	,
(	454	)	,
(	453	)	,
(	453	)	,
(	452	)	,
(	451	)	,
(	450	)	,
(	449	)	,
(	448	)	,
(	447	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	443	)	,
(	442	)	,
(	441	)	,
(	440	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	436	)	,
(	435	)	,
(	434	)	,
(	433	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	429	)	,
(	428	)	,
(	427	)	,
(	426	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	422	)	,
(	421	)	,
(	420	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	416	)	,
(	415	)	,
(	414	)	,
(	413	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	409	)	,
(	408	)	,
(	407	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	403	)	,
(	402	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	398	)	,
(	397	)	,
(	396	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	393	)	,
(	392	)	,
(	391	)	,
(	390	)	,
(	389	)	,
(	389	)	,
(	388	)	,
(	387	)	,
(	386	)	,
(	385	)	,
(	384	)	,
(	384	)	,
(	383	)	,
(	382	)	,
(	381	)	,
(	380	)	,
(	379	)	,
(	379	)	,
(	378	)	,
(	377	)	,
(	376	)	,
(	375	)	,
(	374	)	,
(	374	)	,
(	373	)	,
(	372	)	,
(	371	)	,
(	370	)	,
(	370	)	,
(	369	)	,
(	368	)	,
(	367	)	,
(	366	)	,
(	366	)	,
(	365	)	,
(	364	)	,
(	363	)	,
(	362	)	,
(	361	)	,
(	361	)	,
(	360	)	,
(	359	)	,
(	358	)	,
(	357	)	,
(	357	)	,
(	356	)	,
(	355	)	,
(	354	)	,
(	354	)	,
(	353	)	,
(	352	)	,
(	351	)	,
(	350	)	,
(	350	)	,
(	349	)	,
(	348	)	,
(	347	)	,
(	347	)	,
(	346	)	,
(	345	)	,
(	344	)	,
(	343	)	,
(	343	)	,
(	342	)	,
(	341	)	,
(	340	)	,
(	340	)	,
(	339	)	,
(	338	)	,
(	337	)	,
(	337	)	,
(	336	)	,
(	335	)	,
(	334	)	,
(	334	)	,
(	333	)	,
(	332	)	,
(	331	)	,
(	331	)	,
(	330	)	,
(	329	)	,
(	328	)	,
(	328	)	,
(	327	)	,
(	326	)	,
(	325	)	,
(	325	)	,
(	324	)	,
(	323	)	,
(	323	)	,
(	322	)	,
(	321	)	,
(	320	)	,
(	320	)	,
(	319	)	,
(	318	)	,
(	318	)	,
(	317	)	,
(	316	)	,
(	315	)	,
(	315	)	,
(	314	)	,
(	313	)	,
(	313	)	,
(	312	)	,
(	311	)	,
(	311	)	,
(	310	)	,
(	309	)	,
(	308	)	,
(	308	)	,
(	307	)	,
(	306	)	,
(	306	)	,
(	305	)	,
(	304	)	,
(	304	)	,
(	303	)	,
(	302	)	,
(	302	)	,
(	301	)	,
(	300	)	,
(	300	)	,
(	299	)	,
(	298	)	,
(	298	)	,
(	297	)	,
(	297	)	,
(	296	)	,
(	295	)	,
(	295	)	,
(	294	)	,
(	293	)	,
(	293	)	,
(	292	)	,
(	291	)	,
(	291	)	,
(	290	)	,
(	290	)	,
(	289	)	,
(	288	)	,
(	288	)	,
(	287	)	,
(	286	)	,
(	286	)	,
(	285	)	,
(	285	)	,
(	284	)	,
(	283	)	,
(	283	)	,
(	282	)	,
(	282	)	,
(	281	)	,
(	281	)	,
(	280	)	,
(	279	)	,
(	279	)	,
(	278	)	,
(	278	)	,
(	277	)	,
(	277	)	,
(	276	)	,
(	275	)	,
(	275	)	,
(	274	)	,
(	274	)	,
(	273	)	,
(	273	)	,
(	272	)	,
(	272	)	,
(	271	)	,
(	271	)	,
(	270	)	,
(	269	)	,
(	269	)	,
(	268	)	,
(	268	)	,
(	267	)	,
(	267	)	,
(	266	)	,
(	266	)	,
(	265	)	,
(	265	)	,
(	264	)	,
(	264	)	,
(	263	)	,
(	263	)	,
(	262	)	,
(	262	)	,
(	261	)	,
(	261	)	,
(	260	)	,
(	260	)	,
(	260	)	,
(	259	)	,
(	259	)	,
(	258	)	,
(	258	)	,
(	257	)	,
(	257	)	,
(	256	)	,
(	256	)	,
(	255	)	,
(	255	)	,
(	255	)	,
(	254	)	,
(	254	)	,
(	253	)	,
(	253	)	,
(	252	)	,
(	252	)	,
(	252	)	,
(	251	)	,
(	251	)	,
(	250	)	,
(	250	)	,
(	250	)	,
(	249	)	,
(	249	)	,
(	248	)	,
(	248	)	,
(	248	)	,
(	247	)	,
(	247	)	,
(	247	)	,
(	246	)	,
(	246	)	,
(	245	)	,
(	245	)	,
(	245	)	,
(	244	)	,
(	244	)	,
(	244	)	,
(	243	)	,
(	243	)	,
(	243	)	,
(	242	)	,
(	242	)	,
(	242	)	,
(	242	)	,
(	241	)	,
(	241	)	,
(	241	)	,
(	240	)	,
(	240	)	,
(	240	)	,
(	239	)	,
(	239	)	,
(	239	)	,
(	239	)	,
(	238	)	,
(	238	)	,
(	238	)	,
(	238	)	,
(	237	)	,
(	237	)	,
(	237	)	,
(	237	)	,
(	236	)	,
(	236	)	,
(	236	)	,
(	236	)	,
(	235	)	,
(	235	)	,
(	235	)	,
(	235	)	,
(	235	)	,
(	234	)	,
(	234	)	,
(	234	)	,
(	234	)	,
(	234	)	,
(	233	)	,
(	233	)	,
(	233	)	,
(	233	)	,
(	233	)	,
(	233	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	233	)	,
(	233	)	,
(	233	)	,
(	233	)	,
(	233	)	,
(	234	)	,
(	234	)	,
(	234	)	,
(	234	)	,
(	234	)	,
(	235	)	,
(	235	)	,
(	235	)	,
(	235	)	,
(	236	)	,
(	236	)	,
(	236	)	,
(	236	)	,
(	237	)	,
(	237	)	,
(	237	)	,
(	237	)	,
(	238	)	,
(	238	)	,
(	238	)	,
(	239	)	,
(	239	)	,
(	239	)	,
(	240	)	,
(	240	)	,
(	240	)	,
(	241	)	,
(	241	)	,
(	241	)	,
(	242	)	,
(	242	)	,
(	242	)	,
(	243	)	,
(	243	)	,
(	244	)	,
(	244	)	,
(	244	)	,
(	245	)	,
(	245	)	,
(	246	)	,
(	246	)	,
(	246	)	,
(	247	)	,
(	247	)	,
(	248	)	,
(	248	)	,
(	249	)	,
(	249	)	,
(	250	)	,
(	250	)	,
(	251	)	,
(	251	)	,
(	252	)	,
(	252	)	,
(	253	)	,
(	253	)	,
(	254	)	,
(	254	)	,
(	255	)	,
(	255	)	,
(	256	)	,
(	256	)	,
(	257	)	,
(	258	)	,
(	258	)	,
(	259	)	,
(	259	)	,
(	260	)	,
(	261	)	,
(	261	)	,
(	262	)	,
(	262	)	,
(	263	)	,
(	264	)	,
(	264	)	,
(	265	)	,
(	266	)	,
(	266	)	,
(	267	)	,
(	268	)	,
(	268	)	,
(	269	)	,
(	270	)	,
(	271	)	,
(	271	)	,
(	272	)	,
(	273	)	,
(	273	)	,
(	274	)	,
(	275	)	,
(	276	)	,
(	277	)	,
(	277	)	,
(	278	)	,
(	279	)	,
(	280	)	,
(	280	)	,
(	281	)	,
(	282	)	,
(	283	)	,
(	284	)	,
(	285	)	,
(	285	)	,
(	286	)	,
(	287	)	,
(	288	)	,
(	289	)	,
(	290	)	,
(	291	)	,
(	292	)	,
(	293	)	,
(	293	)	,
(	294	)	,
(	295	)	,
(	296	)	,
(	297	)	,
(	298	)	,
(	299	)	,
(	300	)	,
(	301	)	,
(	302	)	,
(	303	)	,
(	304	)	,
(	305	)	,
(	306	)	,
(	307	)	,
(	308	)	,
(	309	)	,
(	310	)	,
(	311	)	,
(	312	)	,
(	313	)	,
(	314	)	,
(	315	)	,
(	317	)	,
(	318	)	,
(	319	)	,
(	320	)	,
(	321	)	,
(	322	)	,
(	323	)	,
(	324	)	,
(	326	)	,
(	327	)	,
(	328	)	,
(	329	)	,
(	330	)	,
(	332	)	,
(	333	)	,
(	334	)	,
(	335	)	,
(	336	)	,
(	338	)	,
(	339	)	,
(	340	)	,
(	341	)	,
(	343	)	,
(	344	)	,
(	345	)	,
(	347	)	,
(	348	)	,
(	349	)	,
(	351	)	,
(	352	)	,
(	353	)	,
(	355	)	,
(	356	)	,
(	357	)	,
(	359	)	,
(	360	)	,
(	361	)	,
(	363	)	,
(	364	)	,
(	366	)	,
(	367	)	,
(	369	)	,
(	370	)	,
(	371	)	,
(	373	)	,
(	374	)	,
(	376	)	,
(	377	)	,
(	379	)	,
(	380	)	,
(	382	)	,
(	383	)	,
(	385	)	,
(	387	)	,
(	388	)	,
(	390	)	,
(	391	)	,
(	393	)	,
(	394	)	,
(	396	)	,
(	398	)	,
(	399	)	,
(	401	)	,
(	402	)	,
(	404	)	,
(	406	)	,
(	407	)	,
(	409	)	,
(	411	)	,
(	412	)	,
(	414	)	,
(	416	)	,
(	418	)	,
(	419	)	,
(	421	)	,
(	423	)	,
(	425	)	,
(	426	)	,
(	428	)	,
(	430	)	,
(	432	)	,
(	434	)	,
(	435	)	,
(	437	)	,
(	439	)	,
(	441	)	,
(	443	)	,
(	445	)	,
(	447	)	,
(	448	)	,
(	450	)	,
(	452	)	,
(	454	)	,
(	456	)	,
(	458	)	,
(	460	)	,
(	462	)	,
(	464	)	,
(	466	)	,
(	468	)	,
(	470	)	,
(	472	)	,
(	474	)	,
(	476	)	,
(	478	)	,
(	480	)	,
(	482	)	,
(	484	)	,
(	486	)	,
(	488	)	,
(	490	)	,
(	492	)	,
(	495	)	,
(	497	)	,
(	499	)	,
(	501	)	,
(	503	)	,
(	505	)	,
(	508	)	,
(	510	)	,
(	512	)	,
(	514	)	,
(	516	)	,
(	519	)	,
(	521	)	,
(	523	)	,
(	525	)	,
(	528	)	,
(	530	)	,
(	532	)	,
(	535	)	,
(	537	)	,
(	539	)	,
(	542	)	,
(	544	)	,
(	546	)	,
(	549	)	,
(	551	)	,
(	553	)	,
(	556	)	,
(	558	)	,
(	561	)	,
(	563	)	,
(	566	)	,
(	568	)	,
(	570	)	,
(	573	)	,
(	575	)	,
(	578	)	,
(	581	)	,
(	583	)	,
(	586	)	,
(	588	)	,
(	591	)	,
(	593	)	,
(	596	)	,
(	598	)	,
(	601	)	,
(	604	)	,
(	606	)	,
(	609	)	,
(	612	)	,
(	614	)	,
(	617	)	,
(	620	)	,
(	622	)	,
(	625	)	,
(	628	)	,
(	631	)	,
(	633	)	,
(	636	)	,
(	639	)	,
(	642	)	,
(	644	)	,
(	647	)	,
(	650	)	,
(	653	)	,
(	656	)	,
(	659	)	,
(	661	)	,
(	664	)	,
(	667	)	,
(	670	)	,
(	673	)	,
(	676	)	,
(	679	)	,
(	682	)	,
(	685	)	,
(	688	)	,
(	691	)	,
(	694	)	,
(	697	)	,
(	700	)	,
(	703	)	,
(	706	)	,
(	709	)	,
(	712	)	,
(	715	)	,
(	718	)	,
(	721	)	,
(	724	)	,
(	728	)	,
(	731	)	,
(	734	)	,
(	737	)	,
(	740	)	,
(	743	)	,
(	747	)	,
(	750	)	,
(	753	)	,
(	756	)	,
(	760	)	,
(	763	)	,
(	766	)	,
(	770	)	,
(	773	)	,
(	776	)	,
(	780	)	,
(	783	)	,
(	786	)	,
(	790	)	,
(	793	)	,
(	796	)	,
(	800	)	,
(	803	)	,
(	807	)	,
(	810	)	,
(	814	)	,
(	817	)	,
(	821	)	,
(	824	)	,
(	828	)	,
(	831	)	,
(	835	)	,
(	838	)	,
(	842	)	,
(	845	)	,
(	849	)	,
(	853	)	,
(	856	)	,
(	860	)	,
(	864	)	,
(	867	)	,
(	871	)	,
(	875	)	,
(	878	)	,
(	882	)	,
(	886	)	,
(	890	)	,
(	893	)	,
(	897	)	,
(	901	)	,
(	905	)	,
(	909	)	,
(	912	)	,
(	916	)	,
(	920	)	,
(	924	)	,
(	928	)	,
(	932	)	,
(	936	)	,
(	940	)	,
(	944	)	,
(	947	)	,
(	951	)	,
(	955	)	,
(	959	)	,
(	963	)	,
(	967	)	,
(	972	)	,
(	976	)	,
(	980	)	,
(	984	)	,
(	988	)	,
(	992	)	,
(	996	)	,
(	1000	)	,
(	1004	)	,
(	1009	)	,
(	1013	)	,
(	1017	)	,
(	1021	)	,
(	1025	)	,
(	1030	)	,
(	1034	)	,
(	1038	)	,
(	1042	)	,
(	1047	)	,
(	1051	)	,
(	1055	)	,
(	1060	)	,
(	1064	)	,
(	1069	)	,
(	1073	)	,
(	1077	)	,
(	1082	)	,
(	1086	)	,
(	1091	)	,
(	1095	)	,
(	1100	)	,
(	1104	)	,
(	1109	)	,
(	1113	)	,
(	1118	)	,
(	1122	)	,
(	1127	)	,
(	1131	)	,
(	1136	)	,
(	1141	)	,
(	1145	)	,
(	1150	)	,
(	1155	)	,
(	1159	)	,
(	1164	)	,
(	1169	)	,
(	1173	)	,
(	1178	)	,
(	1183	)	,
(	1188	)	,
(	1192	)	,
(	1197	)	,
(	1202	)	,
(	1207	)	,
(	1212	)	,
(	1217	)	,
(	1221	)	,
(	1226	)	,
(	1231	)	,
(	1236	)	,
(	1241	)	,
(	1246	)	,
(	1251	)	,
(	1256	)	,
(	1261	)	,
(	1266	)	,
(	1271	)	,
(	1276	)	,
(	1281	)	,
(	1286	)	,
(	1291	)	,
(	1297	)	,
(	1302	)	,
(	1307	)	,
(	1312	)	,
(	1317	)	,
(	1322	)	,
(	1328	)	,
(	1333	)	,
(	1338	)	,
(	1343	)	,
(	1349	)	,
(	1354	)	,
(	1359	)	,
(	1365	)	,
(	1370	)	,
(	1375	)	,
(	1381	)	,
(	1386	)	,
(	1392	)	,
(	1397	)	,
(	1402	)	,
(	1408	)	,
(	1413	)	,
(	1419	)	,
(	1424	)	,
(	1430	)	,
(	1436	)	,
(	1441	)	,
(	1447	)	,
(	1452	)	,
(	1458	)	,
(	1464	)	,
(	1469	)	,
(	1475	)	,
(	1481	)	,
(	1486	)	,
(	1492	)	,
(	1498	)	,
(	1503	)	,
(	1509	)	,
(	1515	)	,
(	1521	)	,
(	1527	)	,
(	1532	)	,
(	1538	)	,
(	1544	)	,
(	1550	)	,
(	1556	)	,
(	1562	)	,
(	1568	)	,
(	1574	)	,
(	1580	)	,
(	1586	)	,
(	1592	)	,
(	1598	)	,
(	1604	)	,
(	1610	)	,
(	1616	)	,
(	1622	)	,
(	1628	)	,
(	1634	)	,
(	1641	)	,
(	1647	)	,
(	1653	)	,
(	1659	)	,
(	1665	)	,
(	1672	)	,
(	1678	)	,
(	1684	)	,
(	1690	)	,
(	1697	)	,
(	1703	)	,
(	1710	)	,
(	1716	)	,
(	1722	)	,
(	1729	)	,
(	1735	)	,
(	1742	)	,
(	1748	)	,
(	1755	)	,
(	1761	)	,
(	1768	)	,
(	1774	)	,
(	1781	)	,
(	1787	)	,
(	1794	)	,
(	1800	)	,
(	1807	)	,
(	1814	)	,
(	1820	)	,
(	1827	)	,
(	1834	)	,
(	1840	)	,
(	1847	)	,
(	1854	)	,
(	1861	)	,
(	1868	)	,
(	1874	)	,
(	1881	)	,
(	1888	)	,
(	1895	)	,
(	1902	)	,
(	1909	)	,
(	1916	)	,
(	1923	)	,
(	1930	)	,
(	1937	)	,
(	1944	)	,
(	1951	)	,
(	1958	)	,
(	1965	)	,
(	1972	)	,
(	1979	)	,
(	1986	)	,
(	1993	)	,
(	2000	)	,
(	2008	)	,
(	2015	)	,
(	2022	)	,
(	2029	)	,
(	2037	)	,
(	2044	)	,
(	2051	)	,
(	2058	)	,
(	2066	)	,
(	2073	)	,
(	2081	)	,
(	2088	)	,
(	2095	)	,
(	2103	)	,
(	2110	)	,
(	2118	)	,
(	2125	)	,
(	2133	)	,
(	2140	)	,
(	2148	)	,
(	2155	)	,
(	2163	)	,
(	2171	)	,
(	2178	)	,
(	2186	)	,
(	2194	)	,
(	2201	)	,
(	2209	)	,
(	2217	)	,
(	2225	)	,
(	2232	)	,
(	2240	)	,
(	2248	)	,
(	2256	)	,
(	2264	)	,
(	2272	)	,
(	2280	)	,
(	2287	)	,
(	2295	)	,
(	2303	)	,
(	2311	)	,
(	2319	)	,
(	2327	)	,
(	2335	)	,
(	2344	)	,
(	2352	)	,
(	2360	)	,
(	2368	)	,
(	2376	)	,
(	2384	)	,
(	2392	)	,
(	2401	)	,
(	2409	)	,
(	2417	)	,
(	2425	)	,
(	2434	)	,
(	2442	)	,
(	2450	)	,
(	2459	)	,
(	2467	)	,
(	2476	)	,
(	2484	)	,
(	2492	)	,
(	2501	)	,
(	2509	)	,
(	2518	)	,
(	2526	)	,
(	2535	)	,
(	2544	)	,
(	2552	)	,
(	2561	)	,
(	2570	)	,
(	2578	)	,
(	2587	)	,
(	2596	)	,
(	2604	)	,
(	2613	)	,
(	2622	)	,
(	2631	)	,
(	2639	)	,
(	2648	)	,
(	2657	)	,
(	2666	)	,
(	2675	)	,
(	2684	)	,
(	2693	)	,
(	2702	)	,
(	2711	)	,
(	2720	)	,
(	2729	)	,
(	2738	)	,
(	2747	)	,
(	2756	)	,
(	2765	)	,
(	2774	)	,
(	2784	)	,
(	2793	)	,
(	2802	)	,
(	2811	)	,
(	2821	)	,
(	2830	)	,
(	2839	)	,
(	2849	)	,
(	2858	)	,
(	2867	)	,
(	2877	)	,
(	2886	)	,
(	2896	)	,
(	2905	)	,
(	2915	)	,
(	2924	)	,
(	2934	)	,
(	2943	)	,
(	2953	)	,
(	2962	)	,
(	2972	)	,
(	2982	)	,
(	2991	)	,
(	3001	)	,
(	3011	)	,
(	3021	)	,
(	3030	)	,
(	3040	)	,
(	3050	)	,
(	3060	)	,
(	3070	)	,
(	3080	)	,
(	3089	)	,
(	3099	)	,
(	3109	)	,
(	3119	)	,
(	3129	)	,
(	3139	)	,
(	3149	)	,
(	3160	)	,
(	3170	)	,
(	3180	)	,
(	3190	)	,
(	3200	)	,
(	3210	)	,
(	3221	)	,
(	3231	)	,
(	3241	)	,
(	3251	)	,
(	3262	)	,
(	3272	)	,
(	3282	)	,
(	3293	)	,
(	3303	)	,
(	3314	)	,
(	3324	)	,
(	3335	)	,
(	3345	)	,
(	3356	)	,
(	3366	)	,
(	3377	)	,
(	3387	)	,
(	3398	)	,
(	3409	)	,
(	3419	)	,
(	3430	)	,
(	3441	)	,
(	3452	)	,
(	3462	)	,
(	3473	)	,
(	3484	)	,
(	3495	)	,
(	3506	)	,
(	3517	)	,
(	3528	)	,
(	3539	)	,
(	3550	)	,
(	3561	)	,
(	3572	)	,
(	3583	)	,
(	3594	)	,
(	3605	)	,
(	3616	)	,
(	3627	)	,
(	3638	)	,
(	3650	)	,
(	3661	)	,
(	3672	)	,
(	3683	)	,
(	3695	)	,
(	3706	)	,
(	3717	)	,
(	3729	)	,
(	3740	)	,
(	3752	)	,
(	3763	)	,
(	3775	)	,
(	3786	)	,
(	3798	)	,
(	3809	)	,
(	3821	)	,
(	3832	)	,
(	3844	)	,
(	3856	)	,
(	3867	)	,
(	3879	)	,
(	3891	)	,
(	3903	)	,
(	3914	)	,
(	3926	)	,
(	3938	)	,
(	3950	)	,
(	3962	)	,
(	3974	)	,
(	3986	)	,
(	3998	)	,
(	4010	)	,
(	4022	)	,
(	4034	)	,
(	4046	)	,
(	4058	)	,
(	4070	)	,
(	4083	)	,
(	4095	)	,
(	4107	)	,
(	4119	)	,
(	4131	)	,
(	4144	)	,
(	4156	)	,
(	4168	)	,
(	4181	)	,
(	4193	)	,
(	4206	)	,
(	4218	)	,
(	4231	)	,
(	4243	)	,
(	4256	)	,
(	4268	)	,
(	4281	)	,
(	4294	)	,
(	4306	)	,
(	4319	)	,
(	4332	)	,
(	4344	)	,
(	4357	)	,
(	4370	)	,
(	4383	)	,
(	4396	)	,
(	4408	)	,
(	4421	)	,
(	4434	)	,
(	4447	)	,
(	4460	)	,
(	4473	)	,
(	4486	)	,
(	4499	)	,
(	4512	)	,
(	4526	)	,
(	4539	)	,
(	4552	)	,
(	4565	)	,
(	4578	)	,
(	4592	)	,
(	4605	)	,
(	4618	)	,
(	4632	)	,
(	4645	)	,
(	4658	)	,
(	4672	)	,
(	4685	)	,
(	4699	)	,
(	4712	)	,
(	4726	)	,
(	4739	)	,
(	4753	)	,
(	4767	)	,
(	4780	)	,
(	4794	)	,
(	4808	)	,
(	4822	)	,
(	4835	)	,
(	4849	)	,
(	4863	)	,
(	4877	)	,
(	4891	)	,
(	4905	)	,
(	4919	)	,
(	4933	)	,
(	4947	)	,
(	4961	)	,
(	4975	)	,
(	4989	)	,
(	5003	)	,
(	5017	)	,
(	5031	)	,
(	5045	)	,
(	5060	)	,
(	5074	)	,
(	5088	)	,
(	5103	)	,
(	5117	)	,
(	5131	)	,
(	5146	)	,
(	5160	)	,
(	5175	)	,
(	5189	)	,
(	5204	)	,
(	5218	)	,
(	5233	)	,
(	5248	)	,
(	5262	)	,
(	5277	)	,
(	5292	)	,
(	5306	)	,
(	5321	)	,
(	5336	)	,
(	5351	)	,
(	5366	)	,
(	5381	)	,
(	5395	)	,
(	5410	)	,
(	5425	)	,
(	5440	)	,
(	5455	)	,
(	5471	)	,
(	5486	)	,
(	5501	)	,
(	5516	)	,
(	5531	)	,
(	5546	)	,
(	5562	)	,
(	5577	)	,
(	5592	)	,
(	5608	)	,
(	5623	)	,
(	5638	)	,
(	5654	)	,
(	5669	)	,
(	5685	)	,
(	5700	)	,
(	5716	)	,
(	5732	)	,
(	5747	)	,
(	5763	)	,
(	5779	)	,
(	5794	)	,
(	5810	)	,
(	5826	)	,
(	5842	)	,
(	5857	)	,
(	5873	)	,
(	5889	)	,
(	5905	)	,
(	5921	)	,
(	5937	)	,
(	5953	)	,
(	5969	)	,
(	5985	)	,
(	6002	)	,
(	6018	)	,
(	6034	)	,
(	6050	)	,
(	6066	)	,
(	6083	)	,
(	6099	)	,
(	6115	)	,
(	6132	)	,
(	6148	)	,
(	6165	)	,
(	6181	)	,
(	6198	)	,
(	6214	)	,
(	6231	)	,
(	6247	)	,
(	6264	)	,
(	6281	)	,
(	6297	)	,
(	6314	)	,
(	6331	)	,
(	6348	)	,
(	6364	)	,
(	6381	)	,
(	6398	)	,
(	6415	)	,
(	6432	)	,
(	6449	)	,
(	6466	)	,
(	6483	)	,
(	6500	)	,
(	6517	)	,
(	6535	)	,
(	6552	)	,
(	6569	)	,
(	6586	)	,
(	6604	)	,
(	6621	)	,
(	6638	)	,
(	6656	)	,
(	6673	)	,
(	6691	)	,
(	6708	)	,
(	6726	)	,
(	6743	)	,
(	6761	)	,
(	6778	)	,
(	6796	)	,
(	6814	)	,
(	6832	)	,
(	6849	)	,
(	6867	)	,
(	6885	)	,
(	6903	)	,
(	6921	)	,
(	6939	)	,
(	6957	)	,
(	6975	)	,
(	6993	)	,
(	7011	)	,
(	7029	)	,
(	7047	)	,
(	7065	)	,
(	7083	)	,
(	7102	)	,
(	7120	)	,
(	7138	)	,
(	7156	)	,
(	7175	)	,
(	7193	)	,
(	7212	)	,
(	7230	)	,
(	7249	)	,
(	7267	)	,
(	7286	)	,
(	7304	)	,
(	7323	)	,
(	7342	)	,
(	7360	)	,
(	7379	)	,
(	7398	)	,
(	7417	)	,
(	7436	)	,
(	7455	)	,
(	7473	)	,
(	7492	)	,
(	7511	)	,
(	7530	)	,
(	7550	)	,
(	7569	)	,
(	7588	)	,
(	7607	)	,
(	7626	)	,
(	7645	)	,
(	7665	)	,
(	7684	)	,
(	7703	)	,
(	7723	)	,
(	7742	)	,
(	7762	)	,
(	7781	)	,
(	7801	)	,
(	7820	)	,
(	7840	)	,
(	7859	)	,
(	7879	)	,
(	7899	)	,
(	7919	)	,
(	7938	)	,
(	7958	)	,
(	7978	)	,
(	7998	)	,
(	8018	)	,
(	8038	)	,
(	8058	)	,
(	8078	)	,
(	8098	)	,
(	8118	)	,
(	8138	)	,
(	8158	)	,
(	8179	)	,
(	8199	)	,
(	8219	)	,
(	8239	)	,
(	8260	)	,
(	8280	)	,
(	8301	)	,
(	8321	)	,
(	8342	)	,
(	8362	)	,
(	8383	)	,
(	8403	)	,
(	8424	)	,
(	8445	)	,
(	8465	)	,
(	8486	)	,
(	8507	)	,
(	8528	)	,
(	8549	)	,
(	8570	)	,
(	8590	)	,
(	8611	)	,
(	8632	)	,
(	8654	)	,
(	8675	)	,
(	8696	)	,
(	8717	)	,
(	8738	)	,
(	8759	)	,
(	8781	)	,
(	8802	)	,
(	8823	)	,
(	8845	)	,
(	8866	)	,
(	8888	)	,
(	8909	)	,
(	8931	)	,
(	8952	)	,
(	8974	)	,
(	8996	)	,
(	9017	)	,
(	9039	)	,
(	9061	)	,
(	9083	)	,
(	9105	)	,
(	9126	)	,
(	9148	)	,
(	9170	)	,
(	9192	)	,
(	9214	)	,
(	9236	)	,
(	9259	)	,
(	9281	)	,
(	9303	)	,
(	9325	)	,
(	9347	)	,
(	9370	)	,
(	9392	)	,
(	9415	)	,
(	9437	)	,
(	9459	)	,
(	9482	)	,
(	9504	)	,
(	9527	)	,
(	9550	)	,
(	9572	)	,
(	9595	)	,
(	9618	)	,
(	9641	)	,
(	9663	)	,
(	9686	)	,
(	9709	)	,
(	9732	)	,
(	9755	)	,
(	9778	)	,
(	9801	)	,
(	9824	)	,
(	9847	)	,
(	9871	)	,
(	9894	)	,
(	9917	)	,
(	9940	)	,
(	9964	)	,
(	9987	)	,
(	10011	)	,
(	10034	)	,
(	10058	)	,
(	10081	)	,
(	10105	)	,
(	10128	)	,
(	10152	)	,
(	10176	)	,
(	10199	)	,
(	10223	)	,
(	10247	)	,
(	10271	)	,
(	10295	)	,
(	10319	)	,
(	10343	)	,
(	10367	)	,
(	10391	)	,
(	10415	)	,
(	10439	)	,
(	10463	)	,
(	10487	)	,
(	10512	)	,
(	10536	)	,
(	10560	)	,
(	10585	)	,
(	10609	)	,
(	10634	)	,
(	10658	)	,
(	10683	)	,
(	10707	)	,
(	10732	)	,
(	10757	)	,
(	10781	)	,
(	10806	)	,
(	10831	)	,
(	10856	)	,
(	10881	)	,
(	10906	)	,
(	10930	)	,
(	10955	)	,
(	10981	)	,
(	11006	)	,
(	11031	)	,
(	11056	)	,
(	11081	)	,
(	11106	)	,
(	11132	)	,
(	11157	)	,
(	11182	)	,
(	11208	)	,
(	11233	)	,
(	11259	)	,
(	11284	)	,
(	11310	)	,
(	11336	)	,
(	11361	)	,
(	11387	)	,
(	11413	)	,
(	11439	)	,
(	11464	)	,
(	11490	)	,
(	11516	)	,
(	11542	)	,
(	11568	)	,
(	11594	)	,
(	11620	)	,
(	11647	)	,
(	11673	)	,
(	11699	)	,
(	11725	)	,
(	11752	)	,
(	11778	)	,
(	11804	)	,
(	11831	)	,
(	11857	)	,
(	11884	)	,
(	11910	)	,
(	11937	)	,
(	11964	)	,
(	11990	)	,
(	12017	)	,
(	12044	)	,
(	12071	)	,
(	12098	)	,
(	12125	)	,
(	12152	)	,
(	12179	)	,
(	12206	)	,
(	12233	)	,
(	12260	)	,
(	12287	)	,
(	12314	)	,
(	12342	)	,
(	12369	)	,
(	12396	)	,
(	12424	)	,
(	12451	)	,
(	12479	)	,
(	12506	)	,
(	12534	)	,
(	12562	)	,
(	12589	)	,
(	12617	)	,
(	12645	)	,
(	12672	)	,
(	12700	)	,
(	12728	)	,
(	12756	)	,
(	12784	)	,
(	12812	)	,
(	12840	)	,
(	12868	)	,
(	12897	)	,
(	12925	)	,
(	12953	)	,
(	12981	)	,
(	13010	)	,
(	13038	)	,
(	13067	)	,
(	13095	)	,
(	13124	)	,
(	13152	)	,
(	13181	)	,
(	13209	)	,
(	13238	)	,
(	13267	)	,
(	13296	)	,
(	13325	)	,
(	13353	)	,
(	13382	)	,
(	13411	)	,
(	13440	)	,
(	13469	)	,
(	13499	)	,
(	13528	)	,
(	13557	)	,
(	13586	)	,
(	13615	)	,
(	13645	)	,
(	13674	)	,
(	13704	)	,
(	13733	)	,
(	13763	)	,
(	13792	)	,
(	13822	)	,
(	13852	)	,
(	13881	)	,
(	13911	)	,
(	13941	)	,
(	13971	)	,
(	14001	)	,
(	14031	)	,
(	14061	)	,
(	14091	)	,
(	14121	)	,
(	14151	)	,
(	14181	)	,
(	14211	)	,
(	14242	)	,
(	14272	)	,
(	14302	)	,
(	14333	)	,
(	14363	)	,
(	14394	)	,
(	14424	)	,
(	14455	)	,
(	14486	)	,
(	14516	)	,
(	14547	)	,
(	14578	)	,
(	14609	)	,
(	14640	)	,
(	14670	)	,
(	14701	)	,
(	14733	)	,
(	14764	)	,
(	14795	)	,
(	14826	)	,
(	14857	)	,
(	14888	)	,
(	14920	)	,
(	14951	)	,
(	14983	)	,
(	15014	)	,
(	15046	)	,
(	15077	)	,
(	15109	)	,
(	15140	)	,
(	15172	)	,
(	15204	)	,
(	15236	)	,
(	15268	)	,
(	15299	)	,
(	15331	)	,
(	15363	)	,
(	15395	)	,
(	15428	)	,
(	15460	)	,
(	15492	)	,
(	15524	)	,
(	15556	)	,
(	15589	)	,
(	15621	)	,
(	15654	)	,
(	15686	)	,
(	15719	)	,
(	15751	)	,
(	15784	)	,
(	15817	)	,
(	15849	)	,
(	15882	)	,
(	15915	)	,
(	15948	)	,
(	15981	)	,
(	16014	)	,
(	16047	)	,
(	16080	)	,
(	16113	)	,
(	16146	)	,
(	16179	)	,
(	16213	)	,
(	16246	)	,
(	16280	)	,
(	16313	)	,
(	16346	)	,
(	16380	)	,
(	16414	)	,
(	16447	)	,
(	16481	)	,
(	16515	)	,
(	16548	)	,
(	16582	)	,
(	16616	)	,
(	16650	)	,
(	16684	)	,
(	16718	)	,
(	16752	)	,
(	16786	)	,
(	16821	)	,
(	16855	)	,
(	16889	)	,
(	16923	)	,
(	16958	)	,
(	16992	)	,
(	17027	)	,
(	17061	)	,
(	17096	)	,
(	17131	)	,
(	17165	)	,
(	17200	)	,
(	17235	)	,
(	17270	)	,
(	17305	)	,
(	17340	)	,
(	17375	)	,
(	17410	)	,
(	17445	)	,
(	17480	)	,
(	17515	)	,
(	17550	)	,
(	17586	)	,
(	17621	)	,
(	17657	)	,
(	17692	)	,
(	17728	)	,
(	17763	)	,
(	17799	)	,
(	17834	)	,
(	17870	)	,
(	17906	)	,
(	17942	)	,
(	17978	)	,
(	18014	)	,
(	18050	)	,
(	18086	)	,
(	18122	)	,
(	18158	)	,
(	18194	)	,
(	18231	)	,
(	18267	)	,
(	18303	)	,
(	18340	)	,
(	18376	)	,
(	18413	)	,
(	18449	)	,
(	18486	)	,
(	18523	)	,
(	18559	)	,
(	18596	)	,
(	18633	)	,
(	18670	)	,
(	18707	)	,
(	18744	)	,
(	18781	)	,
(	18818	)	,
(	18855	)	,
(	18892	)	,
(	18930	)	,
(	18967	)	,
(	19004	)	,
(	19042	)	,
(	19079	)	,
(	19117	)	,
(	19154	)	,
(	19192	)	,
(	19230	)	,
(	19268	)	,
(	19305	)	,
(	19343	)	,
(	19381	)	,
(	19419	)	,
(	19457	)	,
(	19495	)	,
(	19533	)	,
(	19572	)	,
(	19610	)	,
(	19648	)	,
(	19687	)	,
(	19725	)	,
(	19763	)	,
(	19802	)	,
(	19841	)	,
(	19879	)	,
(	19918	)	,
(	19957	)	,
(	19995	)	,
(	20034	)	,
(	20073	)	,
(	20112	)	,
(	20151	)	,
(	20190	)	,
(	20229	)	,
(	20269	)	,
(	20308	)	,
(	20347	)	,
(	20386	)	,
(	20426	)	,
(	20465	)	,
(	20505	)	,
(	20544	)	,
(	20584	)	,
(	20624	)	,
(	20663	)	,
(	20703	)	,
(	20743	)	,
(	20783	)	,
(	20823	)	,
(	20863	)	,
(	20903	)	,
(	20943	)	,
(	20983	)	,
(	21024	)	,
(	21064	)	,
(	21104	)	,
(	21145	)	,
(	21185	)	,
(	21226	)	,
(	21266	)	,
(	21307	)	,
(	21348	)	,
(	21388	)	,
(	21429	)	,
(	21470	)	,
(	21511	)	,
(	21552	)	,
(	21593	)	,
(	21634	)	,
(	21675	)	,
(	21717	)	,
(	21758	)	,
(	21799	)	,
(	21841	)	,
(	21882	)	,
(	21924	)	,
(	21965	)	,
(	22007	)	,
(	22048	)	,
(	22090	)	,
(	22132	)	,
(	22174	)	,
(	22216	)	,
(	22258	)	,
(	22300	)	,
(	22342	)	,
(	22384	)	,
(	22426	)	,
(	22468	)	,
(	22511	)	,
(	22553	)	,
(	22595	)	,
(	22638	)	,
(	22681	)	,
(	22723	)	,
(	22766	)	,
(	22809	)	,
(	22851	)	,
(	22894	)	,
(	22937	)	,
(	22980	)	,
(	23023	)	,
(	23066	)	,
(	23109	)	,
(	23152	)	,
(	23196	)	,
(	23239	)	,
(	23282	)	,
(	23326	)	,
(	23369	)	,
(	23413	)	,
(	23456	)	,
(	23500	)	,
(	23544	)	,
(	23588	)	,
(	23631	)	,
(	23675	)	,
(	23719	)	,
(	23763	)	,
(	23807	)	,
(	23852	)	,
(	23896	)	,
(	23940	)	,
(	23984	)	,
(	24029	)	,
(	24073	)	,
(	24118	)	,
(	24162	)	,
(	24207	)	,
(	24252	)	,
(	24296	)	,
(	24341	)	,
(	24386	)	,
(	24431	)	,
(	24476	)	,
(	24521	)	,
(	24566	)	,
(	24611	)	,
(	24657	)	,
(	24702	)	,
(	24747	)	,
(	24793	)	,
(	24838	)	,
(	24884	)	,
(	24929	)	,
(	24975	)	,
(	25021	)	,
(	25066	)	,
(	25112	)	,
(	25158	)	,
(	25204	)	,
(	25250	)	,
(	25296	)	,
(	25342	)	,
(	25389	)	,
(	25435	)	,
(	25481	)	,
(	25528	)	,
(	25574	)	,
(	25621	)	,
(	25667	)	,
(	25714	)	,
(	25760	)	,
(	25807	)	,
(	25854	)	,
(	25901	)	,
(	25948	)	,
(	25995	)	,
(	26042	)	,
(	26089	)	,
(	26136	)	,
(	26184	)	,
(	26231	)	,
(	26278	)	,
(	26326	)	,
(	26373	)	,
(	26421	)	,
(	26469	)	,
(	26516	)	,
(	26564	)	,
(	26612	)	,
(	26660	)	,
(	26708	)	,
(	26756	)	,
(	26804	)	,
(	26852	)	,
(	26900	)	,
(	26948	)	,
(	26997	)	,
(	27045	)	,
(	27094	)	,
(	27142	)	,
(	27191	)	,
(	27239	)	,
(	27288	)	,
(	27337	)	,
(	27386	)	,
(	27435	)	,
(	27484	)	,
(	27533	)	,
(	27582	)	,
(	27631	)	,
(	27680	)	,
(	27730	)	,
(	27779	)	,
(	27828	)	,
(	27878	)	,
(	27927	)	,
(	27977	)	,
(	28027	)	,
(	28076	)	,
(	28126	)	,
(	28176	)	,
(	28226	)	,
(	28276	)	,
(	28326	)	,
(	28376	)	,
(	28427	)	,
(	28477	)	,
(	28527	)	,
(	28578	)	,
(	28628	)	,
(	28679	)	,
(	28729	)	,
(	28780	)	,
(	28831	)	,
(	28881	)	,
(	28932	)	,
(	28983	)	,
(	29034	)	,
(	29085	)	,
(	29136	)	,
(	29187	)	,
(	29239	)	,
(	29290	)	,
(	29341	)	,
(	29393	)	,
(	29444	)	,
(	29496	)	,
(	29548	)	,
(	29599	)	,
(	29651	)	,
(	29703	)	,
(	29755	)	,
(	29807	)	,
(	29859	)	,
(	29911	)	,
(	29963	)	,
(	30015	)	,
(	30068	)	,
(	30120	)	,
(	30173	)	,
(	30225	)	,
(	30278	)	,
(	30330	)	,
(	30383	)	,
(	30436	)	,
(	30489	)	,
(	30542	)	,
(	30595	)	,
(	30648	)	,
(	30701	)	,
(	30754	)	,
(	30807	)	,
(	30860	)	,
(	30914	)	,
(	30967	)	,
(	31021	)	,
(	31074	)	,
(	31128	)	,
(	31182	)	,
(	31236	)	,
(	31290	)	,
(	31343	)

);

end package LUT_pkg;
