library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

  (4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4084	)	,
(	4069	)	,
(	4055	)	,
(	4041	)	,
(	4027	)	,
(	4013	)	,
(	3999	)	,
(	3986	)	,
(	3972	)	,
(	3958	)	,
(	3945	)	,
(	3932	)	,
(	3918	)	,
(	3905	)	,
(	3892	)	,
(	3879	)	,
(	3866	)	,
(	3853	)	,
(	3840	)	,
(	3828	)	,
(	3815	)	,
(	3802	)	,
(	3790	)	,
(	3778	)	,
(	3765	)	,
(	3753	)	,
(	3741	)	,
(	3729	)	,
(	3717	)	,
(	3705	)	,
(	3693	)	,
(	3681	)	,
(	3670	)	,
(	3658	)	,
(	3646	)	,
(	3635	)	,
(	3623	)	,
(	3612	)	,
(	3601	)	,
(	3590	)	,
(	3578	)	,
(	3567	)	,
(	3556	)	,
(	3545	)	,
(	3534	)	,
(	3524	)	,
(	3513	)	,
(	3502	)	,
(	3492	)	,
(	3481	)	,
(	3470	)	,
(	3460	)	,
(	3450	)	,
(	3439	)	,
(	3429	)	,
(	3419	)	,
(	3409	)	,
(	3399	)	,
(	3389	)	,
(	3379	)	,
(	3369	)	,
(	3359	)	,
(	3349	)	,
(	3339	)	,
(	3330	)	,
(	3320	)	,
(	3310	)	,
(	3301	)	,
(	3291	)	,
(	3282	)	,
(	3272	)	,
(	3263	)	,
(	3254	)	,
(	3245	)	,
(	3235	)	,
(	3226	)	,
(	3217	)	,
(	3208	)	,
(	3199	)	,
(	3190	)	,
(	3181	)	,
(	3173	)	,
(	3164	)	,
(	3155	)	,
(	3146	)	,
(	3138	)	,
(	3129	)	,
(	3121	)	,
(	3112	)	,
(	3104	)	,
(	3095	)	,
(	3087	)	,
(	3078	)	,
(	3070	)	,
(	3062	)	,
(	3054	)	,
(	3045	)	,
(	3037	)	,
(	3029	)	,
(	3021	)	,
(	3013	)	,
(	3005	)	,
(	2997	)	,
(	2989	)	,
(	2982	)	,
(	2974	)	,
(	2966	)	,
(	2958	)	,
(	2951	)	,
(	2943	)	,
(	2935	)	,
(	2928	)	,
(	2920	)	,
(	2913	)	,
(	2905	)	,
(	2898	)	,
(	2891	)	,
(	2883	)	,
(	2876	)	,
(	2869	)	,
(	2861	)	,
(	2854	)	,
(	2847	)	,
(	2840	)	,
(	2833	)	,
(	2826	)	,
(	2819	)	,
(	2812	)	,
(	2805	)	,
(	2798	)	,
(	2791	)	,
(	2784	)	,
(	2777	)	,
(	2770	)	,
(	2764	)	,
(	2757	)	,
(	2750	)	,
(	2744	)	,
(	2737	)	,
(	2730	)	,
(	2724	)	,
(	2717	)	,
(	2711	)	,
(	2704	)	,
(	2698	)	,
(	2691	)	,
(	2685	)	,
(	2679	)	,
(	2672	)	,
(	2666	)	,
(	2660	)	,
(	2653	)	,
(	2647	)	,
(	2641	)	,
(	2635	)	,
(	2629	)	,
(	2622	)	,
(	2616	)	,
(	2610	)	,
(	2604	)	,
(	2598	)	,
(	2592	)	,
(	2586	)	,
(	2580	)	,
(	2575	)	,
(	2569	)	,
(	2563	)	,
(	2557	)	,
(	2551	)	,
(	2545	)	,
(	2540	)	,
(	2534	)	,
(	2528	)	,
(	2523	)	,
(	2517	)	,
(	2511	)	,
(	2506	)	,
(	2500	)	,
(	2495	)	,
(	2489	)	,
(	2484	)	,
(	2478	)	,
(	2473	)	,
(	2467	)	,
(	2462	)	,
(	2456	)	,
(	2451	)	,
(	2446	)	,
(	2440	)	,
(	2435	)	,
(	2430	)	,
(	2424	)	,
(	2419	)	,
(	2414	)	,
(	2409	)	,
(	2404	)	,
(	2399	)	,
(	2393	)	,
(	2388	)	,
(	2383	)	,
(	2378	)	,
(	2373	)	,
(	2368	)	,
(	2363	)	,
(	2358	)	,
(	2353	)	,
(	2348	)	,
(	2343	)	,
(	2338	)	,
(	2333	)	,
(	2329	)	,
(	2324	)	,
(	2319	)	,
(	2314	)	,
(	2309	)	,
(	2305	)	,
(	2300	)	,
(	2295	)	,
(	2290	)	,
(	2286	)	,
(	2281	)	,
(	2276	)	,
(	2272	)	,
(	2267	)	,
(	2263	)	,
(	2258	)	,
(	2253	)	,
(	2249	)	,
(	2244	)	,
(	2240	)	,
(	2235	)	,
(	2231	)	,
(	2226	)	,
(	2222	)	,
(	2218	)	,
(	2213	)	,
(	2209	)	,
(	2204	)	,
(	2200	)	,
(	2196	)	,
(	2191	)	,
(	2187	)	,
(	2183	)	,
(	2179	)	,
(	2174	)	,
(	2170	)	,
(	2166	)	,
(	2162	)	,
(	2157	)	,
(	2153	)	,
(	2149	)	,
(	2145	)	,
(	2141	)	,
(	2137	)	,
(	2133	)	,
(	2128	)	,
(	2124	)	,
(	2120	)	,
(	2116	)	,
(	2112	)	,
(	2108	)	,
(	2104	)	,
(	2100	)	,
(	2096	)	,
(	2092	)	,
(	2088	)	,
(	2084	)	,
(	2081	)	,
(	2077	)	,
(	2073	)	,
(	2069	)	,
(	2065	)	,
(	2061	)	,
(	2057	)	,
(	2054	)	,
(	2050	)	,
(	2046	)	,
(	2042	)	,
(	2038	)	,
(	2035	)	,
(	2031	)	,
(	2027	)	,
(	2024	)	,
(	2020	)	,
(	2016	)	,
(	2013	)	,
(	2009	)	,
(	2005	)	,
(	2002	)	,
(	1998	)	,
(	1994	)	,
(	1991	)	,
(	1987	)	,
(	1984	)	,
(	1980	)	,
(	1977	)	,
(	1973	)	,
(	1970	)	,
(	1966	)	,
(	1963	)	,
(	1959	)	,
(	1956	)	,
(	1952	)	,
(	1949	)	,
(	1945	)	,
(	1942	)	,
(	1938	)	,
(	1935	)	,
(	1932	)	,
(	1928	)	,
(	1925	)	,
(	1922	)	,
(	1918	)	,
(	1915	)	,
(	1912	)	,
(	1908	)	,
(	1905	)	,
(	1902	)	,
(	1898	)	,
(	1895	)	,
(	1892	)	,
(	1889	)	,
(	1885	)	,
(	1882	)	,
(	1879	)	,
(	1876	)	,
(	1873	)	,
(	1869	)	,
(	1866	)	,
(	1863	)	,
(	1860	)	,
(	1857	)	,
(	1854	)	,
(	1850	)	,
(	1847	)	,
(	1844	)	,
(	1841	)	,
(	1838	)	,
(	1835	)	,
(	1832	)	,
(	1829	)	,
(	1826	)	,
(	1823	)	,
(	1820	)	,
(	1817	)	,
(	1814	)	,
(	1811	)	,
(	1808	)	,
(	1805	)	,
(	1802	)	,
(	1799	)	,
(	1796	)	,
(	1793	)	,
(	1790	)	,
(	1787	)	,
(	1784	)	,
(	1781	)	,
(	1779	)	,
(	1776	)	,
(	1773	)	,
(	1770	)	,
(	1767	)	,
(	1764	)	,
(	1761	)	,
(	1759	)	,
(	1756	)	,
(	1753	)	,
(	1750	)	,
(	1747	)	,
(	1745	)	,
(	1742	)	,
(	1739	)	,
(	1736	)	,
(	1734	)	,
(	1731	)	,
(	1728	)	,
(	1725	)	,
(	1723	)	,
(	1720	)	,
(	1717	)	,
(	1715	)	,
(	1712	)	,
(	1709	)	,
(	1707	)	,
(	1704	)	,
(	1701	)	,
(	1699	)	,
(	1696	)	,
(	1693	)	,
(	1691	)	,
(	1688	)	,
(	1685	)	,
(	1683	)	,
(	1680	)	,
(	1678	)	,
(	1675	)	,
(	1673	)	,
(	1670	)	,
(	1667	)	,
(	1665	)	,
(	1662	)	,
(	1660	)	,
(	1657	)	,
(	1655	)	,
(	1652	)	,
(	1650	)	,
(	1647	)	,
(	1645	)	,
(	1642	)	,
(	1640	)	,
(	1637	)	,
(	1635	)	,
(	1633	)	,
(	1630	)	,
(	1628	)	,
(	1625	)	,
(	1623	)	,
(	1620	)	,
(	1618	)	,
(	1616	)	,
(	1613	)	,
(	1611	)	,
(	1608	)	,
(	1606	)	,
(	1604	)	,
(	1601	)	,
(	1599	)	,
(	1597	)	,
(	1594	)	,
(	1592	)	,
(	1590	)	,
(	1587	)	,
(	1585	)	,
(	1583	)	,
(	1580	)	,
(	1578	)	,
(	1576	)	,
(	1574	)	,
(	1571	)	,
(	1569	)	,
(	1567	)	,
(	1565	)	,
(	1562	)	,
(	1560	)	,
(	1558	)	,
(	1556	)	,
(	1553	)	,
(	1551	)	,
(	1549	)	,
(	1547	)	,
(	1544	)	,
(	1542	)	,
(	1540	)	,
(	1538	)	,
(	1536	)	,
(	1534	)	,
(	1531	)	,
(	1529	)	,
(	1527	)	,
(	1525	)	,
(	1523	)	,
(	1521	)	,
(	1519	)	,
(	1516	)	,
(	1514	)	,
(	1512	)	,
(	1510	)	,
(	1508	)	,
(	1506	)	,
(	1504	)	,
(	1502	)	,
(	1500	)	,
(	1498	)	,
(	1496	)	,
(	1493	)	,
(	1491	)	,
(	1489	)	,
(	1487	)	,
(	1485	)	,
(	1483	)	,
(	1481	)	,
(	1479	)	,
(	1477	)	,
(	1475	)	,
(	1473	)	,
(	1471	)	,
(	1469	)	,
(	1467	)	,
(	1465	)	,
(	1463	)	,
(	1461	)	,
(	1459	)	,
(	1457	)	,
(	1455	)	,
(	1453	)	,
(	1451	)	,
(	1449	)	,
(	1448	)	,
(	1446	)	,
(	1444	)	,
(	1442	)	,
(	1440	)	,
(	1438	)	,
(	1436	)	,
(	1434	)	,
(	1432	)	,
(	1430	)	,
(	1428	)	,
(	1427	)	,
(	1425	)	,
(	1423	)	,
(	1421	)	,
(	1419	)	,
(	1417	)	,
(	1415	)	,
(	1413	)	,
(	1412	)	,
(	1410	)	,
(	1408	)	,
(	1406	)	,
(	1404	)	,
(	1402	)	,
(	1401	)	,
(	1399	)	,
(	1397	)	,
(	1395	)	,
(	1393	)	,
(	1392	)	,
(	1390	)	,
(	1388	)	,
(	1386	)	,
(	1384	)	,
(	1383	)	,
(	1381	)	,
(	1379	)	,
(	1377	)	,
(	1376	)	,
(	1374	)	,
(	1372	)	,
(	1370	)	,
(	1369	)	,
(	1367	)	,
(	1365	)	,
(	1363	)	,
(	1362	)	,
(	1360	)	,
(	1358	)	,
(	1357	)	,
(	1355	)	,
(	1353	)	,
(	1351	)	,
(	1350	)	,
(	1348	)	,
(	1346	)	,
(	1345	)	,
(	1343	)	,
(	1341	)	,
(	1340	)	,
(	1338	)	,
(	1336	)	,
(	1335	)	,
(	1333	)	,
(	1331	)	,
(	1330	)	,
(	1328	)	,
(	1326	)	,
(	1325	)	,
(	1323	)	,
(	1322	)	,
(	1320	)	,
(	1318	)	,
(	1317	)	,
(	1315	)	,
(	1313	)	,
(	1312	)	,
(	1310	)	,
(	1309	)	,
(	1307	)	,
(	1305	)	,
(	1304	)	,
(	1302	)	,
(	1301	)	,
(	1299	)	,
(	1298	)	,
(	1296	)	,
(	1294	)	,
(	1293	)	,
(	1291	)	,
(	1290	)	,
(	1288	)	,
(	1287	)	,
(	1285	)	,
(	1284	)	,
(	1282	)	,
(	1281	)	,
(	1279	)	,
(	1277	)	,
(	1276	)	,
(	1274	)	,
(	1273	)	,
(	1271	)	,
(	1270	)	,
(	1268	)	,
(	1267	)	,
(	1265	)	,
(	1264	)	,
(	1262	)	,
(	1261	)	,
(	1259	)	,
(	1258	)	,
(	1256	)	,
(	1255	)	,
(	1254	)	,
(	1252	)	,
(	1251	)	,
(	1249	)	,
(	1248	)	,
(	1246	)	,
(	1245	)	,
(	1243	)	,
(	1242	)	,
(	1240	)	,
(	1239	)	,
(	1238	)	,
(	1236	)	,
(	1235	)	,
(	1233	)	,
(	1232	)	,
(	1230	)	,
(	1229	)	,
(	1228	)	,
(	1226	)	,
(	1225	)	,
(	1223	)	,
(	1222	)	,
(	1221	)	,
(	1219	)	,
(	1218	)	,
(	1216	)	,
(	1215	)	,
(	1214	)	,
(	1212	)	,
(	1211	)	,
(	1210	)	,
(	1208	)	,
(	1207	)	,
(	1205	)	,
(	1204	)	,
(	1203	)	,
(	1201	)	,
(	1200	)	,
(	1199	)	,
(	1197	)	,
(	1196	)	,
(	1195	)	,
(	1193	)	,
(	1192	)	,
(	1191	)	,
(	1189	)	,
(	1188	)	,
(	1187	)	,
(	1185	)	,
(	1184	)	,
(	1183	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1178	)	,
(	1176	)	,
(	1175	)	,
(	1174	)	,
(	1172	)	,
(	1171	)	,
(	1170	)	,
(	1169	)	,
(	1167	)	,
(	1166	)	,
(	1165	)	,
(	1163	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1158	)	,
(	1157	)	,
(	1156	)	,
(	1155	)	,
(	1153	)	,
(	1152	)	,
(	1151	)	,
(	1150	)	,
(	1148	)	,
(	1147	)	,
(	1146	)	,
(	1145	)	,
(	1143	)	,
(	1142	)	,
(	1141	)	,
(	1140	)	,
(	1139	)	,
(	1137	)	,
(	1136	)	,
(	1135	)	,
(	1134	)	,
(	1132	)	,
(	1131	)	,
(	1130	)	,
(	1129	)	,
(	1128	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1116	)	,
(	1115	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1108	)	,
(	1106	)	,
(	1105	)	,
(	1104	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1098	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1067	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1052	)	,
(	1051	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1025	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1005	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	989	)	,
(	989	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	977	)	,
(	977	)	,
(	976	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	972	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	968	)	,
(	968	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	962	)	,
(	961	)	,
(	961	)	,
(	960	)	,
(	959	)	,
(	958	)	,
(	957	)	,
(	956	)	,
(	955	)	,
(	954	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	951	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	948	)	,
(	947	)	,
(	946	)	,
(	945	)	,
(	944	)	,
(	943	)	,
(	942	)	,
(	942	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	938	)	,
(	937	)	,
(	937	)	,
(	936	)	,
(	935	)	,
(	934	)	,
(	933	)	,
(	932	)	,
(	932	)	,
(	931	)	,
(	930	)	,
(	929	)	,
(	928	)	,
(	927	)	,
(	927	)	,
(	926	)	,
(	925	)	,
(	924	)	,
(	923	)	,
(	923	)	,
(	922	)	,
(	921	)	,
(	920	)	,
(	919	)	,
(	918	)	,
(	918	)	,
(	917	)	,
(	916	)	,
(	915	)	,
(	914	)	,
(	914	)	,
(	913	)	,
(	912	)	,
(	911	)	,
(	910	)	,
(	910	)	,
(	909	)	,
(	908	)	,
(	907	)	,
(	907	)	,
(	906	)	,
(	905	)	,
(	904	)	,
(	903	)	,
(	903	)	,
(	902	)	,
(	901	)	,
(	900	)	,
(	900	)	,
(	899	)	,
(	898	)	,
(	897	)	,
(	896	)	,
(	896	)	,
(	895	)	,
(	894	)	,
(	893	)	,
(	893	)	,
(	892	)	,
(	891	)	,
(	890	)	,
(	890	)	,
(	889	)	,
(	888	)	,
(	887	)	,
(	887	)	,
(	886	)	,
(	885	)	,
(	884	)	,
(	884	)	,
(	883	)	,
(	882	)	,
(	881	)	,
(	881	)	,
(	880	)	,
(	879	)	,
(	878	)	,
(	878	)	,
(	877	)	,
(	876	)	,
(	875	)	,
(	875	)	,
(	874	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	868	)	,
(	867	)	,
(	867	)	,
(	866	)	,
(	865	)	,
(	865	)	,
(	864	)	,
(	863	)	,
(	862	)	,
(	862	)	,
(	861	)	,
(	860	)	,
(	860	)	,
(	859	)	,
(	858	)	,
(	857	)	,
(	857	)	,
(	856	)	,
(	855	)	,
(	855	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	851	)	,
(	850	)	,
(	850	)	,
(	849	)	,
(	848	)	,
(	848	)	,
(	847	)	,
(	846	)	,
(	846	)	,
(	845	)	,
(	844	)	,
(	844	)	,
(	843	)	,
(	842	)	,
(	842	)	,
(	841	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	837	)	,
(	837	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	833	)	,
(	833	)	,
(	832	)	,
(	831	)	,
(	831	)	,
(	830	)	,
(	829	)	,
(	829	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	824	)	,
(	823	)	,
(	822	)	,
(	822	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	816	)	,
(	816	)	,
(	815	)	,
(	814	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	811	)	,
(	811	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	808	)	,
(	807	)	,
(	806	)	,
(	806	)	,
(	805	)	,
(	804	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	796	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	793	)	,
(	793	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	769	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	755	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	747	)	,
(	747	)	,
(	746	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	742	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	729	)	,
(	729	)	,
(	728	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	700	)	,
(	699	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	697	)	,
(	696	)	,
(	696	)	,
(	695	)	,
(	695	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	684	)	,
(	683	)	,
(	683	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	674	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	667	)	,
(	667	)	,
(	666	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	664	)	,
(	664	)	,
(	663	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	661	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	658	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	655	)	,
(	655	)	,
(	654	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	650	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	647	)	,
(	646	)	,
(	646	)	,
(	646	)	,
(	645	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	643	)	,
(	643	)	,
(	642	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	639	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	637	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	635	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	622	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	619	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	617	)	,
(	617	)	,
(	616	)	,
(	616	)	,
(	616	)	,
(	615	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	613	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	610	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	608	)	,
(	607	)	,
(	607	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	601	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	596	)	,
(	596	)	,
(	595	)	,
(	595	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	592	)	,
(	592	)	,
(	591	)	,
(	591	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	586	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	584	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	582	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	579	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	577	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	574	)	,
(	574	)	,
(	574	)	,
(	573	)	,
(	573	)	,
(	573	)	,
(	572	)	,
(	572	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	570	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	567	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	564	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	561	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	559	)	,
(	559	)	,
(	558	)	,
(	558	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	551	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	548	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	539	)	,
(	539	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	537	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	

);

constant d27seg_LUT : array_1d := (
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5000000),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 5555555),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 6250000),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 7142857),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 8333333),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 10000000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 12500000),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 16666666),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 25000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 50000000),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
( 1),
(1)
);

constant d2b_LUT : array_1d := (
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10000 ),
( 10004 ),
( 10006 ),
( 10009 ),
( 10011 ),
( 10014 ),
( 10016 ),
( 10019 ),
( 10021 ),
( 10024 ),
( 10026 ),
( 10029 ),
( 10032 ),
( 10034 ),
( 10037 ),
( 10039 ),
( 10042 ),
( 10044 ),
( 10047 ),
( 10049 ),
( 10052 ),
( 10054 ),
( 10057 ),
( 10060 ),
( 10062 ),
( 10065 ),
( 10067 ),
( 10070 ),
( 10072 ),
( 10075 ),
( 10078 ),
( 10080 ),
( 10083 ),
( 10085 ),
( 10088 ),
( 10090 ),
( 10093 ),
( 10096 ),
( 10098 ),
( 10101 ),
( 10103 ),
( 10106 ),
( 10108 ),
( 10111 ),
( 10114 ),
( 10116 ),
( 10119 ),
( 10121 ),
( 10124 ),
( 10127 ),
( 10129 ),
( 10132 ),
( 10134 ),
( 10137 ),
( 10140 ),
( 10142 ),
( 10145 ),
( 10147 ),
( 10150 ),
( 10153 ),
( 10155 ),
( 10158 ),
( 10160 ),
( 10163 ),
( 10166 ),
( 10168 ),
( 10171 ),
( 10173 ),
( 10176 ),
( 10179 ),
( 10181 ),
( 10184 ),
( 10187 ),
( 10189 ),
( 10192 ),
( 10194 ),
( 10197 ),
( 10200 ),
( 10202 ),
( 10205 ),
( 10208 ),
( 10210 ),
( 10213 ),
( 10215 ),
( 10218 ),
( 10221 ),
( 10223 ),
( 10226 ),
( 10229 ),
( 10231 ),
( 10234 ),
( 10237 ),
( 10239 ),
( 10242 ),
( 10245 ),
( 10247 ),
( 10250 ),
( 10253 ),
( 10255 ),
( 10258 ),
( 10261 ),
( 10263 ),
( 10266 ),
( 10268 ),
( 10271 ),
( 10274 ),
( 10276 ),
( 10279 ),
( 10282 ),
( 10285 ),
( 10287 ),
( 10290 ),
( 10293 ),
( 10295 ),
( 10298 ),
( 10301 ),
( 10303 ),
( 10306 ),
( 10309 ),
( 10311 ),
( 10314 ),
( 10317 ),
( 10319 ),
( 10322 ),
( 10325 ),
( 10327 ),
( 10330 ),
( 10333 ),
( 10336 ),
( 10338 ),
( 10341 ),
( 10344 ),
( 10346 ),
( 10349 ),
( 10352 ),
( 10354 ),
( 10357 ),
( 10360 ),
( 10363 ),
( 10365 ),
( 10368 ),
( 10371 ),
( 10374 ),
( 10376 ),
( 10379 ),
( 10382 ),
( 10384 ),
( 10387 ),
( 10390 ),
( 10393 ),
( 10395 ),
( 10398 ),
( 10401 ),
( 10404 ),
( 10406 ),
( 10409 ),
( 10412 ),
( 10414 ),
( 10417 ),
( 10420 ),
( 10423 ),
( 10425 ),
( 10428 ),
( 10431 ),
( 10434 ),
( 10436 ),
( 10439 ),
( 10442 ),
( 10445 ),
( 10447 ),
( 10450 ),
( 10453 ),
( 10456 ),
( 10459 ),
( 10461 ),
( 10464 ),
( 10467 ),
( 10470 ),
( 10472 ),
( 10475 ),
( 10478 ),
( 10481 ),
( 10483 ),
( 10486 ),
( 10489 ),
( 10492 ),
( 10495 ),
( 10497 ),
( 10500 ),
( 10503 ),
( 10506 ),
( 10509 ),
( 10511 ),
( 10514 ),
( 10517 ),
( 10520 ),
( 10523 ),
( 10525 ),
( 10528 ),
( 10531 ),
( 10534 ),
( 10537 ),
( 10539 ),
( 10542 ),
( 10545 ),
( 10548 ),
( 10551 ),
( 10553 ),
( 10556 ),
( 10559 ),
( 10562 ),
( 10565 ),
( 10567 ),
( 10570 ),
( 10573 ),
( 10576 ),
( 10579 ),
( 10582 ),
( 10584 ),
( 10587 ),
( 10590 ),
( 10593 ),
( 10596 ),
( 10599 ),
( 10601 ),
( 10604 ),
( 10607 ),
( 10610 ),
( 10613 ),
( 10616 ),
( 10619 ),
( 10621 ),
( 10624 ),
( 10627 ),
( 10630 ),
( 10633 ),
( 10636 ),
( 10639 ),
( 10641 ),
( 10644 ),
( 10647 ),
( 10650 ),
( 10653 ),
( 10656 ),
( 10659 ),
( 10661 ),
( 10664 ),
( 10667 ),
( 10670 ),
( 10673 ),
( 10676 ),
( 10679 ),
( 10682 ),
( 10684 ),
( 10687 ),
( 10690 ),
( 10693 ),
( 10696 ),
( 10699 ),
( 10702 ),
( 10705 ),
( 10708 ),
( 10711 ),
( 10713 ),
( 10716 ),
( 10719 ),
( 10722 ),
( 10725 ),
( 10728 ),
( 10731 ),
( 10734 ),
( 10737 ),
( 10740 ),
( 10743 ),
( 10745 ),
( 10748 ),
( 10751 ),
( 10754 ),
( 10757 ),
( 10760 ),
( 10763 ),
( 10766 ),
( 10769 ),
( 10772 ),
( 10775 ),
( 10778 ),
( 10781 ),
( 10784 ),
( 10786 ),
( 10789 ),
( 10792 ),
( 10795 ),
( 10798 ),
( 10801 ),
( 10804 ),
( 10807 ),
( 10810 ),
( 10813 ),
( 10816 ),
( 10819 ),
( 10822 ),
( 10825 ),
( 10828 ),
( 10831 ),
( 10834 ),
( 10837 ),
( 10840 ),
( 10843 ),
( 10846 ),
( 10849 ),
( 10852 ),
( 10855 ),
( 10858 ),
( 10860 ),
( 10863 ),
( 10866 ),
( 10869 ),
( 10872 ),
( 10875 ),
( 10878 ),
( 10881 ),
( 10884 ),
( 10887 ),
( 10890 ),
( 10893 ),
( 10896 ),
( 10899 ),
( 10902 ),
( 10905 ),
( 10908 ),
( 10911 ),
( 10914 ),
( 10917 ),
( 10920 ),
( 10923 ),
( 10926 ),
( 10929 ),
( 10933 ),
( 10936 ),
( 10939 ),
( 10942 ),
( 10945 ),
( 10948 ),
( 10951 ),
( 10954 ),
( 10957 ),
( 10960 ),
( 10963 ),
( 10966 ),
( 10969 ),
( 10972 ),
( 10975 ),
( 10978 ),
( 10981 ),
( 10984 ),
( 10987 ),
( 10990 ),
( 10993 ),
( 10996 ),
( 10999 ),
( 11002 ),
( 11006 ),
( 11009 ),
( 11012 ),
( 11015 ),
( 11018 ),
( 11021 ),
( 11024 ),
( 11027 ),
( 11030 ),
( 11033 ),
( 11036 ),
( 11039 ),
( 11042 ),
( 11045 ),
( 11049 ),
( 11052 ),
( 11055 ),
( 11058 ),
( 11061 ),
( 11064 ),
( 11067 ),
( 11070 ),
( 11073 ),
( 11076 ),
( 11079 ),
( 11083 ),
( 11086 ),
( 11089 ),
( 11092 ),
( 11095 ),
( 11098 ),
( 11101 ),
( 11104 ),
( 11107 ),
( 11111 ),
( 11114 ),
( 11117 ),
( 11120 ),
( 11123 ),
( 11126 ),
( 11129 ),
( 11132 ),
( 11136 ),
( 11139 ),
( 11142 ),
( 11145 ),
( 11148 ),
( 11151 ),
( 11154 ),
( 11158 ),
( 11161 ),
( 11164 ),
( 11167 ),
( 11170 ),
( 11173 ),
( 11177 ),
( 11180 ),
( 11183 ),
( 11186 ),
( 11189 ),
( 11192 ),
( 11195 ),
( 11199 ),
( 11202 ),
( 11205 ),
( 11208 ),
( 11211 ),
( 11215 ),
( 11218 ),
( 11221 ),
( 11224 ),
( 11227 ),
( 11230 ),
( 11234 ),
( 11237 ),
( 11240 ),
( 11243 ),
( 11246 ),
( 11250 ),
( 11253 ),
( 11256 ),
( 11259 ),
( 11262 ),
( 11266 ),
( 11269 ),
( 11272 ),
( 11275 ),
( 11278 ),
( 11282 ),
( 11285 ),
( 11288 ),
( 11291 ),
( 11295 ),
( 11298 ),
( 11301 ),
( 11304 ),
( 11307 ),
( 11311 ),
( 11314 ),
( 11317 ),
( 11320 ),
( 11324 ),
( 11327 ),
( 11330 ),
( 11333 ),
( 11337 ),
( 11340 ),
( 11343 ),
( 11346 ),
( 11350 ),
( 11353 ),
( 11356 ),
( 11359 ),
( 11363 ),
( 11366 ),
( 11369 ),
( 11373 ),
( 11376 ),
( 11379 ),
( 11382 ),
( 11386 ),
( 11389 ),
( 11392 ),
( 11395 ),
( 11399 ),
( 11402 ),
( 11405 ),
( 11409 ),
( 11412 ),
( 11415 ),
( 11418 ),
( 11422 ),
( 11425 ),
( 11428 ),
( 11432 ),
( 11435 ),
( 11438 ),
( 11442 ),
( 11445 ),
( 11448 ),
( 11452 ),
( 11455 ),
( 11458 ),
( 11461 ),
( 11465 ),
( 11468 ),
( 11471 ),
( 11475 ),
( 11478 ),
( 11481 ),
( 11485 ),
( 11488 ),
( 11491 ),
( 11495 ),
( 11498 ),
( 11501 ),
( 11505 ),
( 11508 ),
( 11511 ),
( 11515 ),
( 11518 ),
( 11522 ),
( 11525 ),
( 11528 ),
( 11532 ),
( 11535 ),
( 11538 ),
( 11542 ),
( 11545 ),
( 11548 ),
( 11552 ),
( 11555 ),
( 11559 ),
( 11562 ),
( 11565 ),
( 11569 ),
( 11572 ),
( 11575 ),
( 11579 ),
( 11582 ),
( 11586 ),
( 11589 ),
( 11592 ),
( 11596 ),
( 11599 ),
( 11603 ),
( 11606 ),
( 11609 ),
( 11613 ),
( 11616 ),
( 11620 ),
( 11623 ),
( 11627 ),
( 11630 ),
( 11633 ),
( 11637 ),
( 11640 ),
( 11644 ),
( 11647 ),
( 11650 ),
( 11654 ),
( 11657 ),
( 11661 ),
( 11664 ),
( 11668 ),
( 11671 ),
( 11675 ),
( 11678 ),
( 11681 ),
( 11685 ),
( 11688 ),
( 11692 ),
( 11695 ),
( 11699 ),
( 11702 ),
( 11706 ),
( 11709 ),
( 11713 ),
( 11716 ),
( 11720 ),
( 11723 ),
( 11726 ),
( 11730 ),
( 11733 ),
( 11737 ),
( 11740 ),
( 11744 ),
( 11747 ),
( 11751 ),
( 11754 ),
( 11758 ),
( 11761 ),
( 11765 ),
( 11768 ),
( 11772 ),
( 11775 ),
( 11779 ),
( 11782 ),
( 11786 ),
( 11789 ),
( 11793 ),
( 11796 ),
( 11800 ),
( 11803 ),
( 11807 ),
( 11810 ),
( 11814 ),
( 11818 ),
( 11821 ),
( 11825 ),
( 11828 ),
( 11832 ),
( 11835 ),
( 11839 ),
( 11842 ),
( 11846 ),
( 11849 ),
( 11853 ),
( 11856 ),
( 11860 ),
( 11864 ),
( 11867 ),
( 11871 ),
( 11874 ),
( 11878 ),
( 11881 ),
( 11885 ),
( 11889 ),
( 11892 ),
( 11896 ),
( 11899 ),
( 11903 ),
( 11906 ),
( 11910 ),
( 11914 ),
( 11917 ),
( 11921 ),
( 11924 ),
( 11928 ),
( 11932 ),
( 11935 ),
( 11939 ),
( 11942 ),
( 11946 ),
( 11950 ),
( 11953 ),
( 11957 ),
( 11960 ),
( 11964 ),
( 11968 ),
( 11971 ),
( 11975 ),
( 11979 ),
( 11982 ),
( 11986 ),
( 11989 ),
( 11993 ),
( 11997 ),
( 12000 ),
( 12004 ),
( 12008 ),
( 12011 ),
( 12015 ),
( 12019 ),
( 12022 ),
( 12026 ),
( 12030 ),
( 12033 ),
( 12037 ),
( 12041 ),
( 12044 ),
( 12048 ),
( 12052 ),
( 12055 ),
( 12059 ),
( 12063 ),
( 12066 ),
( 12070 ),
( 12074 ),
( 12077 ),
( 12081 ),
( 12085 ),
( 12088 ),
( 12092 ),
( 12096 ),
( 12099 ),
( 12103 ),
( 12107 ),
( 12111 ),
( 12114 ),
( 12118 ),
( 12122 ),
( 12125 ),
( 12129 ),
( 12133 ),
( 12137 ),
( 12140 ),
( 12144 ),
( 12148 ),
( 12151 ),
( 12155 ),
( 12159 ),
( 12163 ),
( 12166 ),
( 12170 ),
( 12174 ),
( 12178 ),
( 12181 ),
( 12185 ),
( 12189 ),
( 12193 ),
( 12196 ),
( 12200 ),
( 12204 ),
( 12208 ),
( 12212 ),
( 12215 ),
( 12219 ),
( 12223 ),
( 12227 ),
( 12230 ),
( 12234 ),
( 12238 ),
( 12242 ),
( 12246 ),
( 12249 ),
( 12253 ),
( 12257 ),
( 12261 ),
( 12265 ),
( 12268 ),
( 12272 ),
( 12276 ),
( 12280 ),
( 12284 ),
( 12287 ),
( 12291 ),
( 12295 ),
( 12299 ),
( 12303 ),
( 12306 ),
( 12310 ),
( 12314 ),
( 12318 ),
( 12322 ),
( 12326 ),
( 12329 ),
( 12333 ),
( 12337 ),
( 12341 ),
( 12345 ),
( 12349 ),
( 12353 ),
( 12356 ),
( 12360 ),
( 12364 ),
( 12368 ),
( 12372 ),
( 12376 ),
( 12380 ),
( 12384 ),
( 12387 ),
( 12391 ),
( 12395 ),
( 12399 ),
( 12403 ),
( 12407 ),
( 12411 ),
( 12415 ),
( 12419 ),
( 12422 ),
( 12426 ),
( 12430 ),
( 12434 ),
( 12438 ),
( 12442 ),
( 12446 ),
( 12450 ),
( 12454 ),
( 12458 ),
( 12462 ),
( 12465 ),
( 12469 ),
( 12473 ),
( 12477 ),
( 12481 ),
( 12485 ),
( 12489 ),
( 12493 ),
( 12497 ),
( 12501 ),
( 12505 ),
( 12509 ),
( 12513 ),
( 12517 ),
( 12521 ),
( 12525 ),
( 12529 ),
( 12533 ),
( 12537 ),
( 12541 ),
( 12545 ),
( 12548 ),
( 12552 ),
( 12556 ),
( 12560 ),
( 12564 ),
( 12568 ),
( 12572 ),
( 12576 ),
( 12580 ),
( 12584 ),
( 12588 ),
( 12592 ),
( 12596 ),
( 12600 ),
( 12604 ),
( 12608 ),
( 12613 ),
( 12617 ),
( 12621 ),
( 12625 ),
( 12629 ),
( 12633 ),
( 12637 ),
( 12641 ),
( 12645 ),
( 12649 ),
( 12653 ),
( 12657 ),
( 12661 ),
( 12665 ),
( 12669 ),
( 12673 ),
( 12677 ),
( 12681 ),
( 12685 ),
( 12689 ),
( 12693 ),
( 12698 ),
( 12702 ),
( 12706 ),
( 12710 ),
( 12714 ),
( 12718 ),
( 12722 ),
( 12726 ),
( 12730 ),
( 12734 ),
( 12738 ),
( 12743 ),
( 12747 ),
( 12751 ),
( 12755 ),
( 12759 ),
( 12763 ),
( 12767 ),
( 12771 ),
( 12775 ),
( 12780 ),
( 12784 ),
( 12788 ),
( 12792 ),
( 12796 ),
( 12800 ),
( 12804 ),
( 12809 ),
( 12813 ),
( 12817 ),
( 12821 ),
( 12825 ),
( 12829 ),
( 12833 ),
( 12838 ),
( 12842 ),
( 12846 ),
( 12850 ),
( 12854 ),
( 12858 ),
( 12863 ),
( 12867 ),
( 12871 ),
( 12875 ),
( 12879 ),
( 12884 ),
( 12888 ),
( 12892 ),
( 12896 ),
( 12900 ),
( 12905 ),
( 12909 ),
( 12913 ),
( 12917 ),
( 12921 ),
( 12926 ),
( 12930 ),
( 12934 ),
( 12938 ),
( 12943 ),
( 12947 ),
( 12951 ),
( 12955 ),
( 12960 ),
( 12964 ),
( 12968 ),
( 12972 ),
( 12977 ),
( 12981 ),
( 12985 ),
( 12989 ),
( 12994 ),
( 12998 ),
( 13002 ),
( 13006 ),
( 13011 ),
( 13015 ),
( 13019 ),
( 13024 ),
( 13028 ),
( 13032 ),
( 13036 ),
( 13041 ),
( 13045 ),
( 13049 ),
( 13054 ),
( 13058 ),
( 13062 ),
( 13067 ),
( 13071 ),
( 13075 ),
( 13080 ),
( 13084 ),
( 13088 ),
( 13093 ),
( 13097 ),
( 13101 ),
( 13106 ),
( 13110 ),
( 13114 ),
( 13119 ),
( 13123 ),
( 13127 ),
( 13132 ),
( 13136 ),
( 13140 ),
( 13145 ),
( 13149 ),
( 13153 ),
( 13158 ),
( 13162 ),
( 13167 ),
( 13171 ),
( 13175 ),
( 13180 ),
( 13184 ),
( 13189 ),
( 13193 ),
( 13197 ),
( 13202 ),
( 13206 ),
( 13211 ),
( 13215 ),
( 13219 ),
( 13224 ),
( 13228 ),
( 13233 ),
( 13237 ),
( 13242 ),
( 13246 ),
( 13250 ),
( 13255 ),
( 13259 ),
( 13264 ),
( 13268 ),
( 13273 ),
( 13277 ),
( 13282 ),
( 13286 ),
( 13290 ),
( 13295 ),
( 13299 ),
( 13304 ),
( 13308 ),
( 13313 ),
( 13317 ),
( 13322 ),
( 13326 ),
( 13331 ),
( 13335 ),
( 13340 ),
( 13344 ),
( 13349 ),
( 13353 ),
( 13358 ),
( 13362 ),
( 13367 ),
( 13371 ),
( 13376 ),
( 13380 ),
( 13385 ),
( 13389 ),
( 13394 ),
( 13398 ),
( 13403 ),
( 13408 ),
( 13412 ),
( 13417 ),
( 13421 ),
( 13426 ),
( 13430 ),
( 13435 ),
( 13439 ),
( 13444 ),
( 13449 ),
( 13453 ),
( 13458 ),
( 13462 ),
( 13467 ),
( 13471 ),
( 13476 ),
( 13481 ),
( 13485 ),
( 13490 ),
( 13494 ),
( 13499 ),
( 13504 ),
( 13508 ),
( 13513 ),
( 13518 ),
( 13522 ),
( 13527 ),
( 13531 ),
( 13536 ),
( 13541 ),
( 13545 ),
( 13550 ),
( 13555 ),
( 13559 ),
( 13564 ),
( 13569 ),
( 13573 ),
( 13578 ),
( 13582 ),
( 13587 ),
( 13592 ),
( 13597 ),
( 13601 ),
( 13606 ),
( 13611 ),
( 13615 ),
( 13620 ),
( 13625 ),
( 13629 ),
( 13634 ),
( 13639 ),
( 13643 ),
( 13648 ),
( 13653 ),
( 13658 ),
( 13662 ),
( 13667 ),
( 13672 ),
( 13676 ),
( 13681 ),
( 13686 ),
( 13691 ),
( 13695 ),
( 13700 ),
( 13705 ),
( 13710 ),
( 13714 ),
( 13719 ),
( 13724 ),
( 13729 ),
( 13733 ),
( 13738 ),
( 13743 ),
( 13748 ),
( 13752 ),
( 13757 ),
( 13762 ),
( 13767 ),
( 13772 ),
( 13776 ),
( 13781 ),
( 13786 ),
( 13791 ),
( 13796 ),
( 13800 ),
( 13805 ),
( 13810 ),
( 13815 ),
( 13820 ),
( 13825 ),
( 13829 ),
( 13834 ),
( 13839 ),
( 13844 ),
( 13849 ),
( 13854 ),
( 13858 ),
( 13863 ),
( 13868 ),
( 13873 ),
( 13878 ),
( 13883 ),
( 13888 ),
( 13893 ),
( 13897 ),
( 13902 ),
( 13907 ),
( 13912 ),
( 13917 ),
( 13922 ),
( 13927 ),
( 13932 ),
( 13937 ),
( 13941 ),
( 13946 ),
( 13951 ),
( 13956 ),
( 13961 ),
( 13966 ),
( 13971 ),
( 13976 ),
( 13981 ),
( 13986 ),
( 13991 ),
( 13996 ),
( 14001 ),
( 14006 ),
( 14011 ),
( 14016 ),
( 14021 ),
( 14026 ),
( 14030 ),
( 14035 ),
( 14040 ),
( 14045 ),
( 14050 ),
( 14055 ),
( 14060 ),
( 14065 ),
( 14070 ),
( 14075 ),
( 14080 ),
( 14085 ),
( 14090 ),
( 14095 ),
( 14101 ),
( 14106 ),
( 14111 ),
( 14116 ),
( 14121 ),
( 14126 ),
( 14131 ),
( 14136 ),
( 14141 ),
( 14146 ),
( 14151 ),
( 14156 ),
( 14161 ),
( 14166 ),
( 14171 ),
( 14176 ),
( 14181 ),
( 14186 ),
( 14192 ),
( 14197 ),
( 14202 ),
( 14207 ),
( 14212 ),
( 14217 ),
( 14222 ),
( 14227 ),
( 14232 ),
( 14238 ),
( 14243 ),
( 14248 ),
( 14253 ),
( 14258 ),
( 14263 ),
( 14268 ),
( 14273 ),
( 14279 ),
( 14284 ),
( 14289 ),
( 14294 ),
( 14299 ),
( 14304 ),
( 14310 ),
( 14315 ),
( 14320 ),
( 14325 ),
( 14330 ),
( 14336 ),
( 14341 ),
( 14346 ),
( 14351 ),
( 14356 ),
( 14362 ),
( 14367 ),
( 14372 ),
( 14377 ),
( 14382 ),
( 14388 ),
( 14393 ),
( 14398 ),
( 14403 ),
( 14409 ),
( 14414 ),
( 14419 ),
( 14424 ),
( 14430 ),
( 14435 ),
( 14440 ),
( 14445 ),
( 14451 ),
( 14456 ),
( 14461 ),
( 14467 ),
( 14472 ),
( 14477 ),
( 14482 ),
( 14488 ),
( 14493 ),
( 14498 ),
( 14504 ),
( 14509 ),
( 14514 ),
( 14520 ),
( 14525 ),
( 14530 ),
( 14536 ),
( 14541 ),
( 14546 ),
( 14552 ),
( 14557 ),
( 14562 ),
( 14568 ),
( 14573 ),
( 14579 ),
( 14584 ),
( 14589 ),
( 14595 ),
( 14600 ),
( 14605 ),
( 14611 ),
( 14616 ),
( 14622 ),
( 14627 ),
( 14632 ),
( 14638 ),
( 14643 ),
( 14649 ),
( 14654 ),
( 14660 ),
( 14665 ),
( 14670 ),
( 14676 ),
( 14681 ),
( 14687 ),
( 14692 ),
( 14698 ),
( 14703 ),
( 14709 ),
( 14714 ),
( 14720 ),
( 14725 ),
( 14731 ),
( 14736 ),
( 14742 ),
( 14747 ),
( 14753 ),
( 14758 ),
( 14764 ),
( 14769 ),
( 14775 ),
( 14780 ),
( 14786 ),
( 14791 ),
( 14797 ),
( 14802 ),
( 14808 ),
( 14813 ),
( 14819 ),
( 14824 ),
( 14830 ),
( 14836 ),
( 14841 ),
( 14847 ),
( 14852 ),
( 14858 ),
( 14863 ),
( 14869 ),
( 14875 ),
( 14880 ),
( 14886 ),
( 14891 ),
( 14897 ),
( 14903 ),
( 14908 ),
( 14914 ),
( 14919 ),
( 14925 ),
( 14931 ),
( 14936 ),
( 14942 ),
( 14948 ),
( 14953 ),
( 14959 ),
( 14965 ),
( 14970 ),
( 14976 ),
( 14982 ),
( 14987 ),
( 14993 ),
( 14999 ),
( 15004 ),
( 15010 ),
( 15016 ),
( 15021 ),
( 15027 ),
( 15033 ),
( 15039 ),
( 15044 ),
( 15050 ),
( 15056 ),
( 15061 ),
( 15067 ),
( 15073 ),
( 15079 ),
( 15084 ),
( 15090 ),
( 15096 ),
( 15102 ),
( 15107 ),
( 15113 ),
( 15119 ),
( 15125 ),
( 15131 ),
( 15136 ),
( 15142 ),
( 15148 ),
( 15154 ),
( 15160 ),
( 15165 ),
( 15171 ),
( 15177 ),
( 15183 ),
( 15189 ),
( 15194 ),
( 15200 ),
( 15206 ),
( 15212 ),
( 15218 ),
( 15224 ),
( 15230 ),
( 15235 ),
( 15241 ),
( 15247 ),
( 15253 ),
( 15259 ),
( 15265 ),
( 15271 ),
( 15277 ),
( 15283 ),
( 15288 ),
( 15294 ),
( 15300 ),
( 15306 ),
( 15312 ),
( 15318 ),
( 15324 ),
( 15330 ),
( 15336 ),
( 15342 ),
( 15348 ),
( 15354 ),
( 15360 ),
( 15366 ),
( 15372 ),
( 15378 ),
( 15384 ),
( 15390 ),
( 15396 ),
( 15402 ),
( 15408 ),
( 15414 ),
( 15420 ),
( 15426 ),
( 15432 ),
( 15438 ),
( 15444 ),
( 15450 ),
( 15456 ),
( 15462 ),
( 15468 ),
( 15474 ),
( 15480 ),
( 15486 ),
( 15492 ),
( 15498 ),
( 15504 ),
( 15510 ),
( 15516 ),
( 15522 ),
( 15528 ),
( 15535 ),
( 15541 ),
( 15547 ),
( 15553 ),
( 15559 ),
( 15565 ),
( 15571 ),
( 15577 ),
( 15584 ),
( 15590 ),
( 15596 ),
( 15602 ),
( 15608 ),
( 15614 ),
( 15620 ),
( 15627 ),
( 15633 ),
( 15639 ),
( 15645 ),
( 15651 ),
( 15658 ),
( 15664 ),
( 15670 ),
( 15676 ),
( 15682 ),
( 15689 ),
( 15695 ),
( 15701 ),
( 15707 ),
( 15714 ),
( 15720 ),
( 15726 ),
( 15732 ),
( 15739 ),
( 15745 ),
( 15751 ),
( 15757 ),
( 15764 ),
( 15770 ),
( 15776 ),
( 15782 ),
( 15789 ),
( 15795 ),
( 15801 ),
( 15808 ),
( 15814 ),
( 15820 ),
( 15827 ),
( 15833 ),
( 15839 ),
( 15846 ),
( 15852 ),
( 15858 ),
( 15865 ),
( 15871 ),
( 15877 ),
( 15884 ),
( 15890 ),
( 15897 ),
( 15903 ),
( 15909 ),
( 15916 ),
( 15922 ),
( 15929 ),
( 15935 ),
( 15941 ),
( 15948 ),
( 15954 ),
( 15961 ),
( 15967 ),
( 15974 ),
( 15980 ),
( 15987 ),
( 15993 ),
( 16000 ),
( 16006 ),
( 16012 ),
( 16019 ),
( 16025 ),
( 16032 ),
( 16038 ),
( 16045 ),
( 16051 ),
( 16058 ),
( 16064 ),
( 16071 ),
( 16078 ),
( 16084 ),
( 16091 ),
( 16097 ),
( 16104 ),
( 16110 ),
( 16117 ),
( 16123 ),
( 16130 ),
( 16137 ),
( 16143 ),
( 16150 ),
( 16156 ),
( 16163 ),
( 16170 ),
( 16176 ),
( 16183 ),
( 16189 ),
( 16196 ),
( 16203 ),
( 16209 ),
( 16216 ),
( 16223 ),
( 16229 ),
( 16236 ),
( 16243 ),
( 16249 ),
( 16256 ),
( 16263 ),
( 16269 ),
( 16276 ),
( 16283 ),
( 16289 ),
( 16296 ),
( 16303 ),
( 16310 ),
( 16316 ),
( 16323 ),
( 16330 ),
( 16336 ),
( 16343 ),
( 16350 ),
( 16357 ),
( 16363 ),
( 16370 ),
( 16377 ),
( 16384 ),
( 16391 ),
( 16397 ),
( 16404 ),
( 16411 ),
( 16418 ),
( 16425 ),
( 16431 ),
( 16438 ),
( 16445 ),
( 16452 ),
( 16459 ),
( 16466 ),
( 16473 ),
( 16479 ),
( 16486 ),
( 16493 ),
( 16500 ),
( 16507 ),
( 16514 ),
( 16521 ),
( 16528 ),
( 16534 ),
( 16541 ),
( 16548 ),
( 16555 ),
( 16562 ),
( 16569 ),
( 16576 ),
( 16583 ),
( 16590 ),
( 16597 ),
( 16604 ),
( 16611 ),
( 16618 ),
( 16625 ),
( 16632 ),
( 16639 ),
( 16646 ),
( 16653 ),
( 16660 ),
( 16667 ),
( 16674 ),
( 16681 ),
( 16688 ),
( 16695 ),
( 16702 ),
( 16709 ),
( 16716 ),
( 16723 ),
( 16730 ),
( 16737 ),
( 16744 ),
( 16752 ),
( 16759 ),
( 16766 ),
( 16773 ),
( 16780 ),
( 16787 ),
( 16794 ),
( 16801 ),
( 16808 ),
( 16816 ),
( 16823 ),
( 16830 ),
( 16837 ),
( 16844 ),
( 16851 ),
( 16859 ),
( 16866 ),
( 16873 ),
( 16880 ),
( 16887 ),
( 16895 ),
( 16902 ),
( 16909 ),
( 16916 ),
( 16923 ),
( 16931 ),
( 16938 ),
( 16945 ),
( 16953 ),
( 16960 ),
( 16967 ),
( 16974 ),
( 16982 ),
( 16989 ),
( 16996 ),
( 17004 ),
( 17011 ),
( 17018 ),
( 17025 ),
( 17033 ),
( 17040 ),
( 17047 ),
( 17055 ),
( 17062 ),
( 17070 ),
( 17077 ),
( 17084 ),
( 17092 ),
( 17099 ),
( 17106 ),
( 17114 ),
( 17121 ),
( 17129 ),
( 17136 ),
( 17144 ),
( 17151 ),
( 17158 ),
( 17166 ),
( 17173 ),
( 17181 ),
( 17188 ),
( 17196 ),
( 17203 ),
( 17211 ),
( 17218 ),
( 17226 ),
( 17233 ),
( 17241 ),
( 17248 ),
( 17256 ),
( 17263 ),
( 17271 ),
( 17278 ),
( 17286 ),
( 17293 ),
( 17301 ),
( 17309 ),
( 17316 ),
( 17324 ),
( 17331 ),
( 17339 ),
( 17346 ),
( 17354 ),
( 17362 ),
( 17369 ),
( 17377 ),
( 17385 ),
( 17392 ),
( 17400 ),
( 17408 ),
( 17415 ),
( 17423 ),
( 17431 ),
( 17438 ),
( 17446 ),
( 17454 ),
( 17461 ),
( 17469 ),
( 17477 ),
( 17484 ),
( 17492 ),
( 17500 ),
( 17508 ),
( 17515 ),
( 17523 ),
( 17531 ),
( 17539 ),
( 17547 ),
( 17554 ),
( 17562 ),
( 17570 ),
( 17578 ),
( 17586 ),
( 17593 ),
( 17601 ),
( 17609 ),
( 17617 ),
( 17625 ),
( 17633 ),
( 17640 ),
( 17648 ),
( 17656 ),
( 17664 ),
( 17672 ),
( 17680 ),
( 17688 ),
( 17696 ),
( 17704 ),
( 17711 ),
( 17719 ),
( 17727 ),
( 17735 ),
( 17743 ),
( 17751 ),
( 17759 ),
( 17767 ),
( 17775 ),
( 17783 ),
( 17791 ),
( 17799 ),
( 17807 ),
( 17815 ),
( 17823 ),
( 17831 ),
( 17839 ),
( 17847 ),
( 17855 ),
( 17863 ),
( 17872 ),
( 17880 ),
( 17888 ),
( 17896 ),
( 17904 ),
( 17912 ),
( 17920 ),
( 17928 ),
( 17936 ),
( 17944 ),
( 17953 ),
( 17961 ),
( 17969 ),
( 17977 ),
( 17985 ),
( 17993 ),
( 18002 ),
( 18010 ),
( 18018 ),
( 18026 ),
( 18034 ),
( 18043 ),
( 18051 ),
( 18059 ),
( 18067 ),
( 18076 ),
( 18084 ),
( 18092 ),
( 18100 ),
( 18109 ),
( 18117 ),
( 18125 ),
( 18134 ),
( 18142 ),
( 18150 ),
( 18159 ),
( 18167 ),
( 18175 ),
( 18184 ),
( 18192 ),
( 18200 ),
( 18209 ),
( 18217 ),
( 18226 ),
( 18234 ),
( 18242 ),
( 18251 ),
( 18259 ),
( 18268 ),
( 18276 ),
( 18285 ),
( 18293 ),
( 18301 ),
( 18310 ),
( 18318 ),
( 18327 ),
( 18335 ),
( 18344 ),
( 18352 ),
( 18361 ),
( 18369 ),
( 18378 ),
( 18386 ),
( 18395 ),
( 18404 ),
( 18412 ),
( 18421 ),
( 18429 ),
( 18438 ),
( 18446 ),
( 18455 ),
( 18464 ),
( 18472 ),
( 18481 ),
( 18490 ),
( 18498 ),
( 18507 ),
( 18516 ),
( 18524 ),
( 18533 ),
( 18542 ),
( 18550 ),
( 18559 ),
( 18568 ),
( 18576 ),
( 18585 ),
( 18594 ),
( 18603 ),
( 18611 ),
( 18620 ),
( 18629 ),
( 18638 ),
( 18646 ),
( 18655 ),
( 18664 ),
( 18673 ),
( 18682 ),
( 18691 ),
( 18699 ),
( 18708 ),
( 18717 ),
( 18726 ),
( 18735 ),
( 18744 ),
( 18753 ),
( 18761 ),
( 18770 ),
( 18779 ),
( 18788 ),
( 18797 ),
( 18806 ),
( 18815 ),
( 18824 ),
( 18833 ),
( 18842 ),
( 18851 ),
( 18860 ),
( 18869 ),
( 18878 ),
( 18887 ),
( 18896 ),
( 18905 ),
( 18914 ),
( 18923 ),
( 18932 ),
( 18941 ),
( 18950 ),
( 18959 ),
( 18968 ),
( 18977 ),
( 18987 ),
( 18996 ),
( 19005 ),
( 19014 ),
( 19023 ),
( 19032 ),
( 19041 ),
( 19051 ),
( 19060 ),
( 19069 ),
( 19078 ),
( 19087 ),
( 19097 ),
( 19106 ),
( 19115 ),
( 19124 ),
( 19133 ),
( 19143 ),
( 19152 ),
( 19161 ),
( 19171 ),
( 19180 ),
( 19189 ),
( 19198 ),
( 19208 ),
( 19217 ),
( 19226 ),
( 19236 ),
( 19245 ),
( 19255 ),
( 19264 ),
( 19273 ),
( 19283 ),
( 19292 ),
( 19302 ),
( 19311 ),
( 19320 ),
( 19330 ),
( 19339 ),
( 19349 ),
( 19358 ),
( 19368 ),
( 19377 ),
( 19387 ),
( 19396 ),
( 19406 ),
( 19415 ),
( 19425 ),
( 19434 ),
( 19444 ),
( 19453 ),
( 19463 ),
( 19473 ),
( 19482 ),
( 19492 ),
( 19501 ),
( 19511 ),
( 19521 ),
( 19530 ),
( 19540 ),
( 19549 ),
( 19559 ),
( 19569 ),
( 19579 ),
( 19588 ),
( 19598 ),
( 19608 ),
( 19617 ),
( 19627 ),
( 19637 ),
( 19647 ),
( 19656 ),
( 19666 ),
( 19676 ),
( 19686 ),
( 19695 ),
( 19705 ),
( 19715 ),
( 19725 ),
( 19735 ),
( 19745 ),
( 19754 ),
( 19764 ),
( 19774 ),
( 19784 ),
( 19794 ),
( 19804 ),
( 19814 ),
( 19824 ),
( 19834 ),
( 19844 ),
( 19854 ),
( 19864 ),
( 19874 ),
( 19884 ),
( 19894 ),
( 19904 ),
( 19914 ),
( 19924 ),
( 19934 ),
( 19944 ),
( 19954 ),
( 19964 ),
( 19974 ),
( 19984 ),
( 19994 ),
( 20004 ),
( 20014 ),
( 20024 ),
( 20035 ),
( 20045 ),
( 20055 ),
( 20065 ),
( 20075 ),
( 20085 ),
( 20096 ),
( 20106 ),
( 20116 ),
( 20126 ),
( 20137 ),
( 20147 ),
( 20157 ),
( 20167 ),
( 20178 ),
( 20188 ),
( 20198 ),
( 20209 ),
( 20219 ),
( 20229 ),
( 20240 ),
( 20250 ),
( 20260 ),
( 20271 ),
( 20281 ),
( 20292 ),
( 20302 ),
( 20312 ),
( 20323 ),
( 20333 ),
( 20344 ),
( 20354 ),
( 20365 ),
( 20375 ),
( 20386 ),
( 20396 ),
( 20407 ),
( 20417 ),
( 20428 ),
( 20438 ),
( 20449 ),
( 20459 ),
( 20470 ),
( 20481 ),
( 20491 ),
( 20502 ),
( 20512 ),
( 20523 ),
( 20534 ),
( 20544 ),
( 20555 ),
( 20566 ),
( 20576 ),
( 20587 ),
( 20598 ),
( 20609 ),
( 20619 ),
( 20630 ),
( 20641 ),
( 20652 ),
( 20662 ),
( 20673 ),
( 20684 ),
( 20695 ),
( 20706 ),
( 20717 ),
( 20727 ),
( 20738 ),
( 20749 ),
( 20760 ),
( 20771 ),
( 20782 ),
( 20793 ),
( 20804 ),
( 20815 ),
( 20826 ),
( 20837 ),
( 20848 ),
( 20859 ),
( 20870 ),
( 20881 ),
( 20892 ),
( 20903 ),
( 20914 ),
( 20925 ),
( 20936 ),
( 20947 ),
( 20958 ),
( 20969 ),
( 20980 ),
( 20991 ),
( 21003 ),
( 21014 ),
( 21025 ),
( 21036 ),
( 21047 ),
( 21058 ),
( 21070 ),
( 21081 ),
( 21092 ),
( 21103 ),
( 21115 ),
( 21126 ),
( 21137 ),
( 21148 ),
( 21160 ),
( 21171 ),
( 21182 ),
( 21194 ),
( 21205 ),
( 21217 ),
( 21228 ),
( 21239 ),
( 21251 ),
( 21262 ),
( 21274 ),
( 21285 ),
( 21296 ),
( 21308 ),
( 21319 ),
( 21331 ),
( 21342 ),
( 21354 ),
( 21365 ),
( 21377 ),
( 21389 ),
( 21400 ),
( 21412 ),
( 21423 ),
( 21435 ),
( 21447 ),
( 21458 ),
( 21470 ),
( 21482 ),
( 21493 ),
( 21505 ),
( 21517 ),
( 21528 ),
( 21540 ),
( 21552 ),
( 21563 ),
( 21575 ),
( 21587 ),
( 21599 ),
( 21611 ),
( 21622 ),
( 21634 ),
( 21646 ),
( 21658 ),
( 21670 ),
( 21682 ),
( 21694 ),
( 21705 ),
( 21717 ),
( 21729 ),
( 21741 ),
( 21753 ),
( 21765 ),
( 21777 ),
( 21789 ),
( 21801 ),
( 21813 ),
( 21825 ),
( 21837 ),
( 21849 ),
( 21861 ),
( 21873 ),
( 21886 ),
( 21898 ),
( 21910 ),
( 21922 ),
( 21934 ),
( 21946 ),
( 21958 ),
( 21971 ),
( 21983 ),
( 21995 ),
( 22007 ),
( 22020 ),
( 22032 ),
( 22044 ),
( 22056 ),
( 22069 ),
( 22081 ),
( 22093 ),
( 22106 ),
( 22118 ),
( 22130 ),
( 22143 ),
( 22155 ),
( 22168 ),
( 22180 ),
( 22192 ),
( 22205 ),
( 22217 ),
( 22230 ),
( 22242 ),
( 22255 ),
( 22267 ),
( 22280 ),
( 22293 ),
( 22305 ),
( 22318 ),
( 22330 ),
( 22343 ),
( 22356 ),
( 22368 ),
( 22381 ),
( 22393 ),
( 22406 ),
( 22419 ),
( 22432 ),
( 22444 ),
( 22457 ),
( 22470 ),
( 22483 ),
( 22495 ),
( 22508 ),
( 22521 ),
( 22534 ),
( 22547 ),
( 22560 ),
( 22572 ),
( 22585 ),
( 22598 ),
( 22611 ),
( 22624 ),
( 22637 ),
( 22650 ),
( 22663 ),
( 22676 ),
( 22689 ),
( 22702 ),
( 22715 ),
( 22728 ),
( 22741 ),
( 22754 ),
( 22767 ),
( 22780 ),
( 22793 ),
( 22807 ),
( 22820 ),
( 22833 ),
( 22846 ),
( 22859 ),
( 22873 ),
( 22886 ),
( 22899 ),
( 22912 ),
( 22926 ),
( 22939 ),
( 22952 ),
( 22965 ),
( 22979 ),
( 22992 ),
( 23006 ),
( 23019 ),
( 23032 ),
( 23046 ),
( 23059 ),
( 23073 ),
( 23086 ),
( 23100 ),
( 23113 ),
( 23127 ),
( 23140 ),
( 23154 ),
( 23167 ),
( 23181 ),
( 23194 ),
( 23208 ),
( 23222 ),
( 23235 ),
( 23249 ),
( 23263 ),
( 23276 ),
( 23290 ),
( 23304 ),
( 23317 ),
( 23331 ),
( 23345 ),
( 23359 ),
( 23373 ),
( 23386 ),
( 23400 ),
( 23414 ),
( 23428 ),
( 23442 ),
( 23456 ),
( 23470 ),
( 23484 ),
( 23497 ),
( 23511 ),
( 23525 ),
( 23539 ),
( 23553 ),
( 23567 ),
( 23582 ),
( 23596 ),
( 23610 ),
( 23624 ),
( 23638 ),
( 23652 ),
( 23666 ),
( 23680 ),
( 23694 ),
( 23709 ),
( 23723 ),
( 23737 ),
( 23751 ),
( 23766 ),
( 23780 ),
( 23794 ),
( 23809 ),
( 23823 ),
( 23837 ),
( 23852 ),
( 23866 ),
( 23880 ),
( 23895 ),
( 23909 ),
( 23924 ),
( 23938 ),
( 23953 ),
( 23967 ),
( 23982 ),
( 23996 ),
( 24011 ),
( 24025 ),
( 24040 ),
( 24055 ),
( 24069 ),
( 24084 ),
( 24099 ),
( 24113 ),
( 24128 ),
( 24143 ),
( 24158 ),
( 24172 ),
( 24187 ),
( 24202 ),
( 24217 ),
( 24231 ),
( 24246 ),
( 24261 ),
( 24276 ),
( 24291 ),
( 24306 ),
( 24321 ),
( 24336 ),
( 24351 ),
( 24366 ),
( 24381 ),
( 24396 ),
( 24411 ),
( 24426 ),
( 24441 ),
( 24456 ),
( 24471 ),
( 24486 ),
( 24502 ),
( 24517 ),
( 24532 ),
( 24547 ),
( 24562 ),
( 24578 ),
( 24593 ),
( 24608 ),
( 24624 ),
( 24639 ),
( 24654 ),
( 24670 ),
( 24685 ),
( 24701 ),
( 24716 ),
( 24731 ),
( 24747 ),
( 24762 ),
( 24778 ),
( 24793 ),
( 24809 ),
( 24825 ),
( 24840 ),
( 24856 ),
( 24871 ),
( 24887 ),
( 24903 ),
( 24918 ),
( 24934 ),
( 24950 ),
( 24965 ),
( 24981 ),
( 24997 ),
( 25013 ),
( 25029 ),
( 25045 ),
( 25060 ),
( 25076 ),
( 25092 ),
( 25108 ),
( 25124 ),
( 25140 ),
( 25156 ),
( 25172 ),
( 25188 ),
( 25204 ),
( 25220 ),
( 25236 ),
( 25252 ),
( 25268 ),
( 25285 ),
( 25301 ),
( 25317 ),
( 25333 ),
( 25349 ),
( 25366 ),
( 25382 ),
( 25398 ),
( 25415 ),
( 25431 ),
( 25447 ),
( 25464 ),
( 25480 ),
( 25496 ),
( 25513 ),
( 25529 ),
( 25546 ),
( 25562 ),
( 25579 ),
( 25595 ),
( 25612 ),
( 25629 ),
( 25645 ),
( 25662 ),
( 25679 ),
( 25695 ),
( 25712 ),
( 25729 ),
( 25745 ),
( 25762 ),
( 25779 ),
( 25796 ),
( 25813 ),
( 25829 ),
( 25846 ),
( 25863 ),
( 25880 ),
( 25897 ),
( 25914 ),
( 25931 ),
( 25948 ),
( 25965 ),
( 25982 ),
( 25999 ),
( 26016 ),
( 26033 ),
( 26051 ),
( 26068 ),
( 26085 ),
( 26102 ),
( 26119 ),
( 26137 ),
( 26154 ),
( 26171 ),
( 26188 ),
( 26206 ),
( 26223 ),
( 26241 ),
( 26258 ),
( 26275 ),
( 26293 ),
( 26310 ),
( 26328 ),
( 26345 ),
( 26363 ),
( 26381 ),
( 26398 ),
( 26416 ),
( 26433 ),
( 26451 ),
( 26469 ),
( 26487 ),
( 26504 ),
( 26522 ),
( 26540 ),
( 26558 ),
( 26576 ),
( 26593 ),
( 26611 ),
( 26629 ),
( 26647 ),
( 26665 ),
( 26683 ),
( 26701 ),
( 26719 ),
( 26737 ),
( 26755 ),
( 26773 ),
( 26791 ),
( 26810 ),
( 26828 ),
( 26846 ),
( 26864 ),
( 26883 ),
( 26901 ),
( 26919 ),
( 26937 ),
( 26956 ),
( 26974 ),
( 26993 ),
( 27011 ),
( 27029 ),
( 27048 ),
( 27066 ),
( 27085 ),
( 27104 ),
( 27122 ),
( 27141 ),
( 27159 ),
( 27178 ),
( 27197 ),
( 27215 ),
( 27234 ),
( 27253 ),
( 27272 ),
( 27291 ),
( 27309 ),
( 27328 ),
( 27347 ),
( 27366 ),
( 27385 ),
( 27404 ),
( 27423 ),
( 27442 ),
( 27461 ),
( 27480 ),
( 27499 ),
( 27518 ),
( 27537 ),
( 27557 ),
( 27576 ),
( 27595 ),
( 27614 ),
( 27634 ),
( 27653 ),
( 27672 ),
( 27692 ),
( 27711 ),
( 27730 ),
( 27750 ),
( 27769 ),
( 27789 ),
( 27808 ),
( 27828 ),
( 27848 ),
( 27867 ),
( 27887 ),
( 27907 ),
( 27926 ),
( 27946 ),
( 27966 ),
( 27986 ),
( 28005 ),
( 28025 ),
( 28045 ),
( 28065 ),
( 28085 ),
( 28105 ),
( 28125 ),
( 28145 ),
( 28165 ),
( 28185 ),
( 28205 ),
( 28225 ),
( 28245 ),
( 28265 ),
( 28286 ),
( 28306 ),
( 28326 ),
( 28346 ),
( 28367 ),
( 28387 ),
( 28408 ),
( 28428 ),
( 28448 ),
( 28469 ),
( 28489 ),
( 28510 ),
( 28530 ),
( 28551 ),
( 28572 ),
( 28592 ),
( 28613 ),
( 28634 ),
( 28654 ),
( 28675 ),
( 28696 ),
( 28717 ),
( 28738 ),
( 28759 ),
( 28780 ),
( 28800 ),
( 28821 ),
( 28842 ),
( 28863 ),
( 28885 ),
( 28906 ),
( 28927 ),
( 28948 ),
( 28969 ),
( 28990 ),
( 29012 ),
( 29033 ),
( 29054 ),
( 29076 ),
( 29097 ),
( 29118 ),
( 29140 ),
( 29161 ),
( 29183 ),
( 29204 ),
( 29226 ),
( 29248 ),
( 29269 ),
( 29291 ),
( 29313 ),
( 29334 ),
( 29356 ),
( 29378 ),
( 29400 ),
( 29422 ),
( 29444 ),
( 29465 ),
( 29487 ),
( 29509 ),
( 29531 ),
( 29553 ),
( 29576 ),
( 29598 ),
( 29620 ),
( 29642 ),
( 29664 ),
( 29687 ),
( 29709 ),
( 29731 ),
( 29754 ),
( 29776 ),
( 29798 ),
( 29821 ),
( 29843 ),
( 29866 ),
( 29888 ),
( 29911 ),
( 29934 ),
( 29956 ),
( 29979 ),
( 30002 ),
( 30025 ),
( 30047 ),
( 30070 ),
( 30093 ),
( 30116 ),
( 30139 ),
( 30162 ),
( 30185 ),
( 30208 ),
( 30231 ),
( 30254 ),
( 30277 ),
( 30300 ),
( 30324 ),
( 30347 ),
( 30370 ),
( 30394 ),
( 30417 ),
( 30440 ),
( 30464 ),
( 30487 ),
( 30511 ),
( 30534 ),
( 30558 ),
( 30582 ),
( 30605 ),
( 30629 ),
( 30653 ),
( 30676 ),
( 30700 ),
( 30724 ),
( 30748 ),
( 30772 ),
( 30796 ),
( 30820 ),
( 30844 ),
( 30868 ),
( 30892 ),
( 30916 ),
( 30940 ),
( 30965 ),
( 30989 ),
( 31013 ),
( 31037 ),
( 31062 ),
( 31086 ),
( 31111 ),
( 31135 ),
( 31160 ),
( 31184 ),
( 31209 ),
( 31233 ),
( 31258 ),
( 31283 ),
( 31308 ),
( 31332 ),
( 31357 ),
( 31382 ),
( 31407 ),
( 31432 ),
( 31457 ),
( 31482 ),
( 31507 ),
( 31532 ),
( 31557 ),
( 31583 ),
( 31608 ),
( 31633 ),
( 31658 ),
( 31684 ),
( 31709 ),
( 31735 ),
( 31760 ),
( 31786 ),
( 31811 ),
( 31837 ),
( 31862 ),
( 31888 ),
( 31914 ),
( 31940 ),
( 31965 ),
( 31991 ),
( 32017 ),
( 32043 ),
( 32069 ),
( 32095 ),
( 32121 ),
( 32147 ),
( 32173 ),
( 32199 ),
( 32226 ),
( 32252 ),
( 32278 ),
( 32305 ),
( 32331 ),
( 32358 ),
( 32384 ),
( 32411 ),
( 32437 ),
( 32464 ),
( 32490 ),
( 32517 ),
( 32544 ),
( 32571 ),
( 32597 ),
( 32624 ),
( 32651 ),
( 32678 ),
( 32705 ),
( 32732 ),
( 32759 ),
( 32787 ),
( 32814 ),
( 32841 ),
( 32868 ),
( 32896 ),
( 32923 ),
( 32950 ),
( 32978 ),
( 33005 ),
( 33033 ),
( 33061 ),
( 33088 ),
( 33116 ),
( 33144 ),
( 33171 ),
( 33199 ),
( 33227 ),
( 33255 ),
( 33283 ),
( 33311 ),
( 33339 ),
( 33367 ),
( 33395 ),
( 33424 ),
( 33452 ),
( 33480 ),
( 33509 ),
( 33537 ),
( 33565 ),
( 33594 ),
( 33623 ),
( 33651 ),
( 33680 ),
( 33708 ),
( 33737 ),
( 33766 ),
( 33795 ),
( 33824 ),
( 33853 ),
( 33882 ),
( 33911 ),
( 33940 ),
( 33969 ),
( 33998 ),
( 34027 ),
( 34057 ),
( 34086 ),
( 34115 ),
( 34145 ),
( 34174 ),
( 34204 ),
( 34234 ),
( 34263 ),
( 34293 ),
( 34323 ),
( 34352 ),
( 34382 ),
( 34412 ),
( 34442 ),
( 34472 ),
( 34502 ),
( 34532 ),
( 34563 ),
( 34593 ),
( 34623 ),
( 34653 ),
( 34684 ),
( 34714 ),
( 34745 ),
( 34775 ),
( 34806 ),
( 34836 ),
( 34867 ),
( 34898 ),
( 34929 ),
( 34960 ),
( 34991 ),
( 35021 ),
( 35053 ),
( 35084 ),
( 35115 ),
( 35146 ),
( 35177 ),
( 35209 ),
( 35240 ),
( 35271 ),
( 35303 ),
( 35334 ),
( 35366 ),
( 35398 ),
( 35429 ),
( 35461 ),
( 35493 ),
( 35525 ),
( 35557 ),
( 35589 ),
( 35621 ),
( 35653 ),
( 35685 ),
( 35717 ),
( 35749 ),
( 35782 ),
( 35814 ),
( 35847 ),
( 35879 ),
( 35912 ),
( 35944 ),
( 35977 ),
( 36010 ),
( 36043 ),
( 36075 ),
( 36108 ),
( 36141 ),
( 36174 ),
( 36207 ),
( 36241 ),
( 36274 ),
( 36307 ),
( 36341 ),
( 36374 ),
( 36407 ),
( 36441 ),
( 36475 ),
( 36508 ),
( 36542 ),
( 36576 ),
( 36610 ),
( 36643 ),
( 36677 ),
( 36711 ),
( 36746 ),
( 36780 ),
( 36814 ),
( 36848 ),
( 36883 ),
( 36917 ),
( 36952 ),
( 36986 ),
( 37021 ),
( 37055 ),
( 37090 ),
( 37125 ),
( 37160 ),
( 37195 ),
( 37230 ),
( 37265 ),
( 37300 ),
( 37335 ),
( 37370 ),
( 37406 ),
( 37441 ),
( 37477 ),
( 37512 ),
( 37548 ),
( 37583 ),
( 37619 ),
( 37655 ),
( 37691 ),
( 37727 ),
( 37763 ),
( 37799 ),
( 37835 ),
( 37871 ),
( 37908 ),
( 37944 ),
( 37980 ),
( 38017 ),
( 38053 ),
( 38090 ),
( 38127 ),
( 38163 ),
( 38200 ),
( 38237 ),
( 38274 ),
( 38311 ),
( 38348 ),
( 38386 ),
( 38423 ),
( 38460 ),
( 38498 ),
( 38535 ),
( 38573 ),
( 38610 ),
( 38648 ),
( 38686 ),
( 38724 ),
( 38762 ),
( 38800 ),
( 38838 ),
( 38876 ),
( 38914 ),
( 38953 ),
( 38991 ),
( 39029 ),
( 39068 ),
( 39107 ),
( 39145 ),
( 39184 ),
( 39223 ),
( 39262 ),
( 39301 ),
( 39340 ),
( 39379 ),
( 39418 ),
( 39458 ),
( 39497 ),
( 39537 ),
( 39576 ),
( 39616 ),
( 39655 ),
( 39695 ),
( 39735 ),
( 39775 ),
( 39815 ),
( 39855 ),
( 39895 ),
( 39936 ),
( 39976 ),
( 40016 ),
( 40057 ),
( 40098 ),
( 40138 ),
( 40179 ),
( 40220 ),
( 40261 ),
( 40302 ),
( 40343 ),
( 40384 ),
( 40425 ),
( 40467 ),
( 40508 ),
( 40550 ),
( 40591 ),
( 40633 ),
( 40675 ),
( 40717 ),
( 40759 ),
( 40801 ),
( 40843 ),
( 40885 ),
( 40927 ),
( 40970 ),
( 41012 ),
( 41055 ),
( 41097 ),
( 41140 ),
( 41183 ),
( 41226 ),
( 41269 ),
( 41312 ),
( 41355 ),
( 41398 ),
( 41442 ),
( 41485 ),
( 41529 ),
( 41572 ),
( 41616 ),
( 41660 ),
( 41704 ),
( 41748 ),
( 41792 ),
( 41836 ),
( 41880 ),
( 41925 ),
( 41969 ),
( 42014 ),
( 42059 ),
( 42103 ),
( 42148 ),
( 42193 ),
( 42238 ),
( 42283 ),
( 42329 ),
( 42374 ),
( 42419 ),
( 42465 ),
( 42510 ),
( 42556 ),
( 42602 ),
( 42648 ),
( 42694 ),
( 42740 ),
( 42786 ),
( 42833 ),
( 42879 ),
( 42926 ),
( 42972 ),
( 43019 ),
( 43066 ),
( 43113 ),
( 43160 ),
( 43207 ),
( 43254 ),
( 43301 ),
( 43349 ),
( 43396 ),
( 43444 ),
( 43492 ),
( 43540 ),
( 43588 ),
( 43636 ),
( 43684 ),
( 43732 ),
( 43781 ),
( 43829 ),
( 43878 ),
( 43927 ),
( 43975 ),
( 44024 ),
( 44073 ),
( 44123 ),
( 44172 ),
( 44221 ),
( 44271 ),
( 44320 ),
( 44370 ),
( 44420 ),
( 44470 ),
( 44520 ),
( 44570 ),
( 44620 ),
( 44671 ),
( 44721 ),
( 44772 ),
( 44822 ),
( 44873 ),
( 44924 ),
( 44975 ),
( 45026 ),
( 45078 ),
( 45129 ),
( 45181 ),
( 45232 ),
( 45284 ),
( 45336 ),
( 45388 ),
( 45440 ),
( 45492 ),
( 45545 ),
( 45597 ),
( 45650 ),
( 45703 ),
( 45756 ),
( 45809 ),
( 45862 ),
( 45915 ),
( 45968 ),
( 46022 ),
( 46075 ),
( 46129 ),
( 46183 ),
( 46237 ),
( 46291 ),
( 46345 ),
( 46400 ),
( 46454 ),
( 46509 ),
( 46563 ),
( 46618 ),
( 46673 ),
( 46728 ),
( 46784 ),
( 46839 ),
( 46895 ),
( 46950 ),
( 47006 ),
( 47062 ),
( 47118 ),
( 47174 ),
( 47230 ),
( 47287 ),
( 47344 ),
( 47400 ),
( 47457 ),
( 47514 ),
( 47571 ),
( 47628 ),
( 47686 ),
( 47743 ),
( 47801 ),
( 47859 ),
( 47917 ),
( 47975 ),
( 48033 ),
( 48092 ),
( 48150 ),
( 48209 ),
( 48268 ),
( 48327 ),
( 48386 ),
( 48445 ),
( 48504 ),
( 48564 ),
( 48624 ),
( 48684 ),
( 48744 ),
( 48804 ),
( 48864 ),
( 48924 ),
( 48985 ),
( 49046 ),
( 49107 ),
( 49168 ),
( 49229 ),
( 49290 ),
( 49352 ),
( 49413 ),
( 49475 ),
( 49537 ),
( 49599 ),
( 49661 ),
( 49724 ),
( 49786 ),
( 49849 ),
( 49912 ),
( 49975 ),
( 50038 ),
( 50102 ),
( 50165 ),
( 50229 ),
( 50293 ),
( 50357 ),
( 50421 ),
( 50485 ),
( 50550 ),
( 50614 ),
( 50679 ),
( 50744 ),
( 50809 ),
( 50875 ),
( 50940 ),
( 51006 ),
( 51072 ),
( 51138 ),
( 51204 ),
( 51270 ),
( 51337 ),
( 51404 ),
( 51470 ),
( 51538 ),
( 51605 ),
( 51672 ),
( 51740 ),
( 51808 ),
( 51875 ),
( 51944 ),
( 52012 ),
( 52080 ),
( 52149 ),
( 52218 ),
( 52287 ),
( 52356 ),
( 52425 ),
( 52495 ),
( 52565 ),
( 52635 ),
( 52705 ),
( 52775 ),
( 52846 ),
( 52916 ),
( 52987 ),
( 53058 ),
( 53129 ),
( 53201 ),
( 53273 ),
( 53344 ),
( 53416 ),
( 53489 ),
( 53561 ),
( 53634 ),
( 53706 ),
( 53780 ),
( 53853 ),
( 53926 ),
( 54000 ),
( 54074 ),
( 54148 ),
( 54222 ),
( 54296 ),
( 54371 ),
( 54446 ),
( 54521 ),
( 54596 ),
( 54671 ),
( 54747 ),
( 54823 ),
( 54899 ),
( 54975 ),
( 55052 ),
( 55128 ),
( 55205 ),
( 55283 ),
( 55360 ),
( 55437 ),
( 55515 ),
( 55593 ),
( 55672 ),
( 55750 ),
( 55829 ),
( 55908 ),
( 55987 ),
( 56066 ),
( 56146 ),
( 56225 ),
( 56305 ),
( 56386 ),
( 56466 ),
( 56547 ),
( 56628 ),
( 56709 ),
( 56790 ),
( 56872 ),
( 56954 ),
( 57036 ),
( 57118 ),
( 57201 ),
( 57284 ),
( 57367 ),
( 57450 ),
( 57534 ),
( 57618 ),
( 57702 ),
( 57786 ),
( 57870 ),
( 57955 ),
( 58040 ),
( 58125 ),
( 58211 ),
( 58297 ),
( 58383 ),
( 58469 ),
( 58556 ),
( 58642 ),
( 58729 ),
( 58817 ),
( 58904 ),
( 58992 ),
( 59080 ),
( 59169 ),
( 59257 ),
( 59346 ),
( 59435 ),
( 59525 ),
( 59614 ),
( 59704 ),
( 59795 ),
( 59885 ),
( 59976 ),
( 60067 ),
( 60158 ),
( 60250 ),
( 60342 ),
( 60434 ),
( 60527 ),
( 60619 ),
( 60712 ),
( 60806 ),
( 60899 ),
( 60993 ),
( 61087 ),
( 61182 ),
( 61277 ),
( 61372 ),
( 61467 ),
( 61563 ),
( 61659 ),
( 61755 ),
( 61851 ),
( 61948 ),
( 62045 ),
( 62143 ),
( 62241 ),
( 62339 ),
( 62437 ),
( 62536 ),
( 62635 ),
( 62734 ),
( 62834 ),
( 62934 ),
( 63034 ),
( 63135 ),
( 63236 ),
( 63337 ),
( 63438 ),
( 63540 ),
( 63642 ),
( 63745 ),
( 63848 ),
( 63951 ),
( 64055 ),
( 64159 ),
( 64263 ),
( 64367 ),
( 64472 ),
( 64577 ),
( 64683 ),
( 64789 ),
( 64895 ),
( 65002 ),
( 65109 ),
( 65216 ),
( 65324 ),
( 65432 ),
( 65540 ),
( 65649 ),
( 65758 ),
( 65868 ),
( 65978 ),
( 66088 ),
( 66198 ),
( 66309 ),
( 66421 ),
( 66532 ),
( 66644 ),
( 66757 ),
( 66870 ),
( 66983 ),
( 67097 ),
( 67211 ),
( 67325 ),
( 67440 ),
( 67555 ),
( 67670 ),
( 67786 ),
( 67903 ),
( 68019 ),
( 68137 ),
( 68254 ),
( 68372 ),
( 68491 ),
( 68609 ),
( 68729 ),
( 68848 ),
( 68968 ),
( 69089 ),
( 69209 ),
( 69331 ),
( 69452 ),
( 69575 ),
( 69697 ),
( 69820 ),
( 69944 ),
( 70068 ),
( 70192 ),
( 70317 ),
( 70442 ),
( 70567 ),
( 70694 ),
( 70820 ),
( 70947 ),
( 71075 ),
( 71203 ),
( 71331 ),
( 71460 ),
( 71589 ),
( 71719 ),
( 71849 ),
( 71980 ),
( 72111 ),
( 72243 ),
( 72375 ),
( 72508 ),
( 72641 ),
( 72774 ),
( 72908 ),
( 73043 ),
( 73178 ),
( 73314 ),
( 73450 ),
( 73587 ),
( 73724 ),
( 73861 ),
( 73999 ),
( 74138 ),
( 74277 ),
( 74417 ),
( 74557 ),
( 74698 ),
( 74839 ),
( 74981 ),
( 75124 ),
( 75267 ),
( 75410 ),
( 75554 ),
( 75699 ),
( 75844 ),
( 75989 ),
( 76136 ),
( 76282 ),
( 76430 ),
( 76578 ),
( 76726 ),
( 76875 ),
( 77025 ),
( 77175 ),
( 77326 ),
( 77478 ),
( 77630 ),
( 77782 ),
( 77936 ),
( 78089 ),
( 78244 ),
( 78399 ),
( 78555 ),
( 78711 ),
( 78868 ),
( 79025 ),
( 79184 ),
( 79342 ),
( 79502 ),
( 79662 ),
( 79823 ),
( 79984 ),
( 80146 ),
( 80309 ),
( 80472 ),
( 80636 ),
( 80801 ),
( 80966 ),
( 81132 ),
( 81299 ),
( 81466 ),
( 81635 ),
( 81803 ),
( 81973 ),
( 82143 ),
( 82314 ),
( 82486 ),
( 82658 ),
( 82831 ),
( 83005 ),
( 83179 ),
( 83355 ),
( 83531 ),
( 83707 ),
( 83885 ),
( 84063 ),
( 84242 ),
( 84422 ),
( 84602 ),
( 84784 ),
( 84966 ),
( 85149 ),
( 85332 ),
( 85517 ),
( 85702 ),
( 85888 ),
( 86075 ),
( 86263 ),
( 86451 ),
( 86641 ),
( 86831 ),
( 87022 ),
( 87214 ),
( 87406 ),
( 87600 ),
( 87794 ),
( 87989 ),
( 88186 ),
( 88383 ),
( 88580 ),
( 88779 ),
( 88979 ),
( 89180 ),
( 89381 ),
( 89583 ),
( 89787 ),
( 89991 ),
( 90196 ),
( 90402 ),
( 90609 ),
( 90817 ),
( 91026 ),
( 91236 ),
( 91447 ),
( 91659 ),
( 91872 ),
( 92086 ),
( 92301 ),
( 92516 ),
( 92733 ),
( 92951 ),
( 93170 ),
( 93390 ),
( 93611 ),
( 93833 ),
( 94056 ),
( 94280 ),
( 94506 ),
( 94732 ),
( 94959 ),
( 95188 ),
( 95417 ),
( 95648 ),
( 95880 ),
( 96113 ),
( 96347 ),
( 96582 ),
( 96818 ),
( 97056 ),
( 97295 ),
( 97535 ),
( 97776 ),
( 98018 ),
( 98261 ),
( 98506 ),
( 98752 ),
( 98999 ),
( 99247 ),
( 99497 ),
( 99748 ),
( 100000 ),
( 100253 ),
( 100508 ),
( 100764 ),
( 101021 ),
( 101280 ),
( 101540 ),
( 101801 ),
( 102064 ),
( 102328 ),
( 102593 ),
( 102860 ),
( 103128 ),
( 103398 ),
( 103669 ),
( 103941 ),
( 104215 ),
( 104490 ),
( 104767 ),
( 105045 ),
( 105325 ),
( 105606 ),
( 105889 ),
( 106173 ),
( 106458 ),
( 106746 ),
( 107035 ),
( 107325 ),
( 107617 ),
( 107910 ),
( 108206 ),
( 108502 ),
( 108801 ),
( 109101 ),
( 109403 ),
( 109706 ),
( 110011 ),
( 110318 ),
( 110626 ),
( 110936 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 ),
( 166666 )
);




end package LUT_pkg;
