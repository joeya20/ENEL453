library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (
(	6745	)	,
(	6731	)	,
(	6718	)	,
(	6704	)	,
(	6690	)	,
(	6677	)	,
(	6663	)	,
(	6650	)	,
(	6637	)	,
(	6623	)	,
(	6610	)	,
(	6596	)	,
(	6583	)	,
(	6570	)	,
(	6556	)	,
(	6543	)	,
(	6530	)	,
(	6517	)	,
(	6504	)	,
(	6490	)	,
(	6477	)	,
(	6464	)	,
(	6451	)	,
(	6438	)	,
(	6425	)	,
(	6412	)	,
(	6399	)	,
(	6386	)	,
(	6373	)	,
(	6360	)	,
(	6347	)	,
(	6334	)	,
(	6321	)	,
(	6309	)	,
(	6296	)	,
(	6283	)	,
(	6270	)	,
(	6258	)	,
(	6245	)	,
(	6232	)	,
(	6219	)	,
(	6207	)	,
(	6194	)	,
(	6182	)	,
(	6169	)	,
(	6156	)	,
(	6144	)	,
(	6131	)	,
(	6119	)	,
(	6106	)	,
(	6094	)	,
(	6082	)	,
(	6069	)	,
(	6057	)	,
(	6045	)	,
(	6032	)	,
(	6020	)	,
(	6008	)	,
(	5995	)	,
(	5983	)	,
(	5971	)	,
(	5959	)	,
(	5947	)	,
(	5934	)	,
(	5922	)	,
(	5910	)	,
(	5898	)	,
(	5886	)	,
(	5874	)	,
(	5862	)	,
(	5850	)	,
(	5838	)	,
(	5826	)	,
(	5814	)	,
(	5802	)	,
(	5791	)	,
(	5779	)	,
(	5767	)	,
(	5755	)	,
(	5743	)	,
(	5732	)	,
(	5720	)	,
(	5708	)	,
(	5696	)	,
(	5685	)	,
(	5673	)	,
(	5662	)	,
(	5650	)	,
(	5638	)	,
(	5627	)	,
(	5615	)	,
(	5604	)	,
(	5592	)	,
(	5581	)	,
(	5569	)	,
(	5558	)	,
(	5547	)	,
(	5535	)	,
(	5524	)	,
(	5512	)	,
(	5501	)	,
(	5490	)	,
(	5479	)	,
(	5467	)	,
(	5456	)	,
(	5445	)	,
(	5434	)	,
(	5423	)	,
(	5411	)	,
(	5400	)	,
(	5389	)	,
(	5378	)	,
(	5367	)	,
(	5356	)	,
(	5345	)	,
(	5334	)	,
(	5323	)	,
(	5312	)	,
(	5301	)	,
(	5290	)	,
(	5279	)	,
(	5269	)	,
(	5258	)	,
(	5247	)	,
(	5236	)	,
(	5225	)	,
(	5215	)	,
(	5204	)	,
(	5193	)	,
(	5182	)	,
(	5172	)	,
(	5161	)	,
(	5150	)	,
(	5140	)	,
(	5129	)	,
(	5119	)	,
(	5108	)	,
(	5098	)	,
(	5087	)	,
(	5077	)	,
(	5066	)	,
(	5056	)	,
(	5045	)	,
(	5035	)	,
(	5024	)	,
(	5014	)	,
(	5004	)	,
(	4993	)	,
(	4983	)	,
(	4973	)	,
(	4962	)	,
(	4952	)	,
(	4942	)	,
(	4932	)	,
(	4922	)	,
(	4911	)	,
(	4901	)	,
(	4891	)	,
(	4881	)	,
(	4871	)	,
(	4861	)	,
(	4851	)	,
(	4841	)	,
(	4831	)	,
(	4821	)	,
(	4811	)	,
(	4801	)	,
(	4791	)	,
(	4781	)	,
(	4771	)	,
(	4761	)	,
(	4752	)	,
(	4742	)	,
(	4732	)	,
(	4722	)	,
(	4712	)	,
(	4703	)	,
(	4693	)	,
(	4683	)	,
(	4673	)	,
(	4664	)	,
(	4654	)	,
(	4645	)	,
(	4635	)	,
(	4625	)	,
(	4616	)	,
(	4606	)	,
(	4597	)	,
(	4587	)	,
(	4578	)	,
(	4568	)	,
(	4559	)	,
(	4549	)	,
(	4540	)	,
(	4530	)	,
(	4521	)	,
(	4512	)	,
(	4502	)	,
(	4493	)	,
(	4484	)	,
(	4474	)	,
(	4465	)	,
(	4456	)	,
(	4447	)	,
(	4438	)	,
(	4428	)	,
(	4419	)	,
(	4410	)	,
(	4401	)	,
(	4392	)	,
(	4383	)	,
(	4374	)	,
(	4364	)	,
(	4355	)	,
(	4346	)	,
(	4337	)	,
(	4328	)	,
(	4319	)	,
(	4311	)	,
(	4302	)	,
(	4293	)	,
(	4284	)	,
(	4275	)	,
(	4266	)	,
(	4257	)	,
(	4248	)	,
(	4240	)	,
(	4231	)	,
(	4222	)	,
(	4213	)	,
(	4205	)	,
(	4196	)	,
(	4187	)	,
(	4178	)	,
(	4170	)	,
(	4161	)	,
(	4153	)	,
(	4144	)	,
(	4135	)	,
(	4127	)	,
(	4118	)	,
(	4110	)	,
(	4101	)	,
(	4093	)	,
(	4084	)	,
(	4076	)	,
(	4067	)	,
(	4059	)	,
(	4050	)	,
(	4042	)	,
(	4034	)	,
(	4025	)	,
(	4017	)	,
(	4009	)	,
(	4000	)	,
(	3992	)	,
(	3984	)	,
(	3976	)	,
(	3967	)	,
(	3959	)	,
(	3951	)	,
(	3943	)	,
(	3935	)	,
(	3926	)	,
(	3918	)	,
(	3910	)	,
(	3902	)	,
(	3894	)	,
(	3886	)	,
(	3878	)	,
(	3870	)	,
(	3862	)	,
(	3854	)	,
(	3846	)	,
(	3838	)	,
(	3830	)	,
(	3822	)	,
(	3814	)	,
(	3806	)	,
(	3798	)	,
(	3791	)	,
(	3783	)	,
(	3775	)	,
(	3767	)	,
(	3759	)	,
(	3751	)	,
(	3744	)	,
(	3736	)	,
(	3728	)	,
(	3721	)	,
(	3713	)	,
(	3705	)	,
(	3698	)	,
(	3690	)	,
(	3682	)	,
(	3675	)	,
(	3667	)	,
(	3659	)	,
(	3652	)	,
(	3644	)	,
(	3637	)	,
(	3629	)	,
(	3622	)	,
(	3614	)	,
(	3607	)	,
(	3599	)	,
(	3592	)	,
(	3585	)	,
(	3577	)	,
(	3570	)	,
(	3563	)	,
(	3555	)	,
(	3548	)	,
(	3541	)	,
(	3533	)	,
(	3526	)	,
(	3519	)	,
(	3511	)	,
(	3504	)	,
(	3497	)	,
(	3490	)	,
(	3483	)	,
(	3475	)	,
(	3468	)	,
(	3461	)	,
(	3454	)	,
(	3447	)	,
(	3440	)	,
(	3433	)	,
(	3426	)	,
(	3419	)	,
(	3412	)	,
(	3405	)	,
(	3398	)	,
(	3391	)	,
(	3384	)	,
(	3377	)	,
(	3370	)	,
(	3363	)	,
(	3356	)	,
(	3349	)	,
(	3342	)	,
(	3335	)	,
(	3328	)	,
(	3322	)	,
(	3315	)	,
(	3308	)	,
(	3301	)	,
(	3294	)	,
(	3288	)	,
(	3281	)	,
(	3274	)	,
(	3267	)	,
(	3261	)	,
(	3254	)	,
(	3247	)	,
(	3241	)	,
(	3234	)	,
(	3227	)	,
(	3221	)	,
(	3214	)	,
(	3208	)	,
(	3201	)	,
(	3195	)	,
(	3188	)	,
(	3182	)	,
(	3175	)	,
(	3169	)	,
(	3162	)	,
(	3156	)	,
(	3149	)	,
(	3143	)	,
(	3136	)	,
(	3130	)	,
(	3124	)	,
(	3117	)	,
(	3111	)	,
(	3104	)	,
(	3098	)	,
(	3092	)	,
(	3086	)	,
(	3079	)	,
(	3073	)	,
(	3067	)	,
(	3060	)	,
(	3054	)	,
(	3048	)	,
(	3042	)	,
(	3036	)	,
(	3030	)	,
(	3023	)	,
(	3017	)	,
(	3011	)	,
(	3005	)	,
(	2999	)	,
(	2993	)	,
(	2987	)	,
(	2981	)	,
(	2975	)	,
(	2969	)	,
(	2963	)	,
(	2957	)	,
(	2951	)	,
(	2945	)	,
(	2939	)	,
(	2933	)	,
(	2927	)	,
(	2921	)	,
(	2915	)	,
(	2909	)	,
(	2903	)	,
(	2897	)	,
(	2891	)	,
(	2886	)	,
(	2880	)	,
(	2874	)	,
(	2868	)	,
(	2862	)	,
(	2857	)	,
(	2851	)	,
(	2845	)	,
(	2839	)	,
(	2834	)	,
(	2828	)	,
(	2822	)	,
(	2817	)	,
(	2811	)	,
(	2805	)	,
(	2800	)	,
(	2794	)	,
(	2788	)	,
(	2783	)	,
(	2777	)	,
(	2772	)	,
(	2766	)	,
(	2761	)	,
(	2755	)	,
(	2750	)	,
(	2744	)	,
(	2739	)	,
(	2733	)	,
(	2728	)	,
(	2722	)	,
(	2717	)	,
(	2711	)	,
(	2706	)	,
(	2701	)	,
(	2695	)	,
(	2690	)	,
(	2684	)	,
(	2679	)	,
(	2674	)	,
(	2668	)	,
(	2663	)	,
(	2658	)	,
(	2653	)	,
(	2647	)	,
(	2642	)	,
(	2637	)	,
(	2632	)	,
(	2626	)	,
(	2621	)	,
(	2616	)	,
(	2611	)	,
(	2606	)	,
(	2600	)	,
(	2595	)	,
(	2590	)	,
(	2585	)	,
(	2580	)	,
(	2575	)	,
(	2570	)	,
(	2565	)	,
(	2560	)	,
(	2555	)	,
(	2550	)	,
(	2544	)	,
(	2539	)	,
(	2534	)	,
(	2530	)	,
(	2525	)	,
(	2520	)	,
(	2515	)	,
(	2510	)	,
(	2505	)	,
(	2500	)	,
(	2495	)	,
(	2490	)	,
(	2485	)	,
(	2480	)	,
(	2475	)	,
(	2471	)	,
(	2466	)	,
(	2461	)	,
(	2456	)	,
(	2451	)	,
(	2447	)	,
(	2442	)	,
(	2437	)	,
(	2432	)	,
(	2428	)	,
(	2423	)	,
(	2418	)	,
(	2413	)	,
(	2409	)	,
(	2404	)	,
(	2399	)	,
(	2395	)	,
(	2390	)	,
(	2386	)	,
(	2381	)	,
(	2376	)	,
(	2372	)	,
(	2367	)	,
(	2363	)	,
(	2358	)	,
(	2353	)	,
(	2349	)	,
(	2344	)	,
(	2340	)	,
(	2335	)	,
(	2331	)	,
(	2326	)	,
(	2322	)	,
(	2317	)	,
(	2313	)	,
(	2309	)	,
(	2304	)	,
(	2300	)	,
(	2295	)	,
(	2291	)	,
(	2287	)	,
(	2282	)	,
(	2278	)	,
(	2273	)	,
(	2269	)	,
(	2265	)	,
(	2260	)	,
(	2256	)	,
(	2252	)	,
(	2248	)	,
(	2243	)	,
(	2239	)	,
(	2235	)	,
(	2231	)	,
(	2226	)	,
(	2222	)	,
(	2218	)	,
(	2214	)	,
(	2210	)	,
(	2205	)	,
(	2201	)	,
(	2197	)	,
(	2193	)	,
(	2189	)	,
(	2185	)	,
(	2181	)	,
(	2176	)	,
(	2172	)	,
(	2168	)	,
(	2164	)	,
(	2160	)	,
(	2156	)	,
(	2152	)	,
(	2148	)	,
(	2144	)	,
(	2140	)	,
(	2136	)	,
(	2132	)	,
(	2128	)	,
(	2124	)	,
(	2120	)	,
(	2116	)	,
(	2112	)	,
(	2108	)	,
(	2104	)	,
(	2101	)	,
(	2097	)	,
(	2093	)	,
(	2089	)	,
(	2085	)	,
(	2081	)	,
(	2077	)	,
(	2073	)	,
(	2070	)	,
(	2066	)	,
(	2062	)	,
(	2058	)	,
(	2054	)	,
(	2051	)	,
(	2047	)	,
(	2043	)	,
(	2039	)	,
(	2036	)	,
(	2032	)	,
(	2028	)	,
(	2025	)	,
(	2021	)	,
(	2017	)	,
(	2013	)	,
(	2010	)	,
(	2006	)	,
(	2002	)	,
(	1999	)	,
(	1995	)	,
(	1992	)	,
(	1988	)	,
(	1984	)	,
(	1981	)	,
(	1977	)	,
(	1974	)	,
(	1970	)	,
(	1967	)	,
(	1963	)	,
(	1959	)	,
(	1956	)	,
(	1952	)	,
(	1949	)	,
(	1945	)	,
(	1942	)	,
(	1938	)	,
(	1935	)	,
(	1932	)	,
(	1928	)	,
(	1925	)	,
(	1921	)	,
(	1918	)	,
(	1914	)	,
(	1911	)	,
(	1908	)	,
(	1904	)	,
(	1901	)	,
(	1897	)	,
(	1894	)	,
(	1891	)	,
(	1887	)	,
(	1884	)	,
(	1881	)	,
(	1877	)	,
(	1874	)	,
(	1871	)	,
(	1868	)	,
(	1864	)	,
(	1861	)	,
(	1858	)	,
(	1855	)	,
(	1851	)	,
(	1848	)	,
(	1845	)	,
(	1842	)	,
(	1838	)	,
(	1835	)	,
(	1832	)	,
(	1829	)	,
(	1826	)	,
(	1823	)	,
(	1819	)	,
(	1816	)	,
(	1813	)	,
(	1810	)	,
(	1807	)	,
(	1804	)	,
(	1801	)	,
(	1798	)	,
(	1794	)	,
(	1791	)	,
(	1788	)	,
(	1785	)	,
(	1782	)	,
(	1779	)	,
(	1776	)	,
(	1773	)	,
(	1770	)	,
(	1767	)	,
(	1764	)	,
(	1761	)	,
(	1758	)	,
(	1755	)	,
(	1752	)	,
(	1749	)	,
(	1746	)	,
(	1743	)	,
(	1740	)	,
(	1737	)	,
(	1735	)	,
(	1732	)	,
(	1729	)	,
(	1726	)	,
(	1723	)	,
(	1720	)	,
(	1717	)	,
(	1714	)	,
(	1711	)	,
(	1709	)	,
(	1706	)	,
(	1703	)	,
(	1700	)	,
(	1697	)	,
(	1694	)	,
(	1692	)	,
(	1689	)	,
(	1686	)	,
(	1683	)	,
(	1681	)	,
(	1678	)	,
(	1675	)	,
(	1672	)	,
(	1670	)	,
(	1667	)	,
(	1664	)	,
(	1661	)	,
(	1659	)	,
(	1656	)	,
(	1653	)	,
(	1651	)	,
(	1648	)	,
(	1645	)	,
(	1643	)	,
(	1640	)	,
(	1637	)	,
(	1635	)	,
(	1632	)	,
(	1629	)	,
(	1627	)	,
(	1624	)	,
(	1622	)	,
(	1619	)	,
(	1616	)	,
(	1614	)	,
(	1611	)	,
(	1609	)	,
(	1606	)	,
(	1604	)	,
(	1601	)	,
(	1599	)	,
(	1596	)	,
(	1593	)	,
(	1591	)	,
(	1588	)	,
(	1586	)	,
(	1583	)	,
(	1581	)	,
(	1579	)	,
(	1576	)	,
(	1574	)	,
(	1571	)	,
(	1569	)	,
(	1566	)	,
(	1564	)	,
(	1561	)	,
(	1559	)	,
(	1557	)	,
(	1554	)	,
(	1552	)	,
(	1549	)	,
(	1547	)	,
(	1545	)	,
(	1542	)	,
(	1540	)	,
(	1537	)	,
(	1535	)	,
(	1533	)	,
(	1530	)	,
(	1528	)	,
(	1526	)	,
(	1523	)	,
(	1521	)	,
(	1519	)	,
(	1517	)	,
(	1514	)	,
(	1512	)	,
(	1510	)	,
(	1507	)	,
(	1505	)	,
(	1503	)	,
(	1501	)	,
(	1498	)	,
(	1496	)	,
(	1494	)	,
(	1492	)	,
(	1490	)	,
(	1487	)	,
(	1485	)	,
(	1483	)	,
(	1481	)	,
(	1479	)	,
(	1476	)	,
(	1474	)	,
(	1472	)	,
(	1470	)	,
(	1468	)	,
(	1466	)	,
(	1463	)	,
(	1461	)	,
(	1459	)	,
(	1457	)	,
(	1455	)	,
(	1453	)	,
(	1451	)	,
(	1449	)	,
(	1446	)	,
(	1444	)	,
(	1442	)	,
(	1440	)	,
(	1438	)	,
(	1436	)	,
(	1434	)	,
(	1432	)	,
(	1430	)	,
(	1428	)	,
(	1426	)	,
(	1424	)	,
(	1422	)	,
(	1420	)	,
(	1418	)	,
(	1416	)	,
(	1414	)	,
(	1412	)	,
(	1410	)	,
(	1408	)	,
(	1406	)	,
(	1404	)	,
(	1402	)	,
(	1400	)	,
(	1398	)	,
(	1396	)	,
(	1394	)	,
(	1392	)	,
(	1390	)	,
(	1388	)	,
(	1387	)	,
(	1385	)	,
(	1383	)	,
(	1381	)	,
(	1379	)	,
(	1377	)	,
(	1375	)	,
(	1373	)	,
(	1371	)	,
(	1370	)	,
(	1368	)	,
(	1366	)	,
(	1364	)	,
(	1362	)	,
(	1360	)	,
(	1358	)	,
(	1357	)	,
(	1355	)	,
(	1353	)	,
(	1351	)	,
(	1349	)	,
(	1348	)	,
(	1346	)	,
(	1344	)	,
(	1342	)	,
(	1340	)	,
(	1339	)	,
(	1337	)	,
(	1335	)	,
(	1333	)	,
(	1332	)	,
(	1330	)	,
(	1328	)	,
(	1326	)	,
(	1325	)	,
(	1323	)	,
(	1321	)	,
(	1320	)	,
(	1318	)	,
(	1316	)	,
(	1314	)	,
(	1313	)	,
(	1311	)	,
(	1309	)	,
(	1308	)	,
(	1306	)	,
(	1304	)	,
(	1303	)	,
(	1301	)	,
(	1299	)	,
(	1298	)	,
(	1296	)	,
(	1295	)	,
(	1293	)	,
(	1291	)	,
(	1290	)	,
(	1288	)	,
(	1286	)	,
(	1285	)	,
(	1283	)	,
(	1282	)	,
(	1280	)	,
(	1278	)	,
(	1277	)	,
(	1275	)	,
(	1274	)	,
(	1272	)	,
(	1271	)	,
(	1269	)	,
(	1267	)	,
(	1266	)	,
(	1264	)	,
(	1263	)	,
(	1261	)	,
(	1260	)	,
(	1258	)	,
(	1257	)	,
(	1255	)	,
(	1254	)	,
(	1252	)	,
(	1251	)	,
(	1249	)	,
(	1248	)	,
(	1246	)	,
(	1245	)	,
(	1243	)	,
(	1242	)	,
(	1240	)	,
(	1239	)	,
(	1237	)	,
(	1236	)	,
(	1234	)	,
(	1233	)	,
(	1232	)	,
(	1230	)	,
(	1229	)	,
(	1227	)	,
(	1226	)	,
(	1224	)	,
(	1223	)	,
(	1222	)	,
(	1220	)	,
(	1219	)	,
(	1217	)	,
(	1216	)	,
(	1215	)	,
(	1213	)	,
(	1212	)	,
(	1210	)	,
(	1209	)	,
(	1208	)	,
(	1206	)	,
(	1205	)	,
(	1204	)	,
(	1202	)	,
(	1201	)	,
(	1199	)	,
(	1198	)	,
(	1197	)	,
(	1195	)	,
(	1194	)	,
(	1193	)	,
(	1191	)	,
(	1190	)	,
(	1189	)	,
(	1188	)	,
(	1186	)	,
(	1185	)	,
(	1184	)	,
(	1182	)	,
(	1181	)	,
(	1180	)	,
(	1178	)	,
(	1177	)	,
(	1176	)	,
(	1175	)	,
(	1173	)	,
(	1172	)	,
(	1171	)	,
(	1170	)	,
(	1168	)	,
(	1167	)	,
(	1166	)	,
(	1165	)	,
(	1163	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1158	)	,
(	1157	)	,
(	1156	)	,
(	1155	)	,
(	1154	)	,
(	1152	)	,
(	1151	)	,
(	1150	)	,
(	1149	)	,
(	1148	)	,
(	1146	)	,
(	1145	)	,
(	1144	)	,
(	1143	)	,
(	1142	)	,
(	1141	)	,
(	1139	)	,
(	1138	)	,
(	1137	)	,
(	1136	)	,
(	1135	)	,
(	1134	)	,
(	1132	)	,
(	1131	)	,
(	1130	)	,
(	1129	)	,
(	1128	)	,
(	1127	)	,
(	1126	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1121	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1116	)	,
(	1115	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1105	)	,
(	1104	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1099	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1090	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1080	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1069	)	,
(	1068	)	,
(	1067	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1054	)	,
(	1053	)	,
(	1052	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1045	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1031	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1025	)	,
(	1025	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1020	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1016	)	,
(	1016	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1012	)	,
(	1012	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1005	)	,
(	1004	)	,
(	1004	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	1000	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	994	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	991	)	,
(	990	)	,
(	989	)	,
(	988	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	985	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	979	)	,
(	979	)	,
(	978	)	,
(	977	)	,
(	977	)	,
(	976	)	,
(	975	)	,
(	974	)	,
(	974	)	,
(	973	)	,
(	972	)	,
(	972	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	969	)	,
(	968	)	,
(	967	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	962	)	,
(	962	)	,
(	961	)	,
(	960	)	,
(	960	)	,
(	959	)	,
(	958	)	,
(	958	)	,
(	957	)	,
(	956	)	,
(	956	)	,
(	955	)	,
(	954	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	952	)	,
(	951	)	,
(	950	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	948	)	,
(	947	)	,
(	946	)	,
(	946	)	,
(	945	)	,
(	944	)	,
(	944	)	,
(	943	)	,
(	942	)	,
(	942	)	,
(	941	)	,
(	940	)	,
(	940	)	,
(	939	)	,
(	939	)	,
(	938	)	,
(	937	)	,
(	937	)	,
(	936	)	,
(	935	)	,
(	935	)	,
(	934	)	,
(	933	)	,
(	933	)	,
(	932	)	,
(	932	)	,
(	931	)	,
(	930	)	,
(	930	)	,
(	929	)	,
(	928	)	,
(	928	)	,
(	927	)	,
(	927	)	,
(	926	)	,
(	925	)	,
(	925	)	,
(	924	)	,
(	923	)	,
(	923	)	,
(	922	)	,
(	922	)	,
(	921	)	,
(	920	)	,
(	920	)	,
(	919	)	,
(	919	)	,
(	918	)	,
(	917	)	,
(	917	)	,
(	916	)	,
(	915	)	,
(	915	)	,
(	914	)	,
(	914	)	,
(	913	)	,
(	912	)	,
(	912	)	,
(	911	)	,
(	911	)	,
(	910	)	,
(	909	)	,
(	909	)	,
(	908	)	,
(	908	)	,
(	907	)	,
(	907	)	,
(	906	)	,
(	905	)	,
(	905	)	,
(	904	)	,
(	904	)	,
(	903	)	,
(	902	)	,
(	902	)	,
(	901	)	,
(	901	)	,
(	900	)	,
(	899	)	,
(	899	)	,
(	898	)	,
(	898	)	,
(	897	)	,
(	897	)	,
(	896	)	,
(	895	)	,
(	895	)	,
(	894	)	,
(	894	)	,
(	893	)	,
(	893	)	,
(	892	)	,
(	891	)	,
(	891	)	,
(	890	)	,
(	890	)	,
(	889	)	,
(	888	)	,
(	888	)	,
(	887	)	,
(	887	)	,
(	886	)	,
(	886	)	,
(	885	)	,
(	885	)	,
(	884	)	,
(	883	)	,
(	883	)	,
(	882	)	,
(	882	)	,
(	881	)	,
(	881	)	,
(	880	)	,
(	879	)	,
(	879	)	,
(	878	)	,
(	878	)	,
(	877	)	,
(	877	)	,
(	876	)	,
(	875	)	,
(	875	)	,
(	874	)	,
(	874	)	,
(	873	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	869	)	,
(	868	)	,
(	868	)	,
(	867	)	,
(	867	)	,
(	866	)	,
(	865	)	,
(	865	)	,
(	864	)	,
(	864	)	,
(	863	)	,
(	863	)	,
(	862	)	,
(	862	)	,
(	861	)	,
(	860	)	,
(	860	)	,
(	859	)	,
(	859	)	,
(	858	)	,
(	858	)	,
(	857	)	,
(	857	)	,
(	856	)	,
(	856	)	,
(	855	)	,
(	854	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	852	)	,
(	851	)	,
(	851	)	,
(	850	)	,
(	850	)	,
(	849	)	,
(	848	)	,
(	848	)	,
(	847	)	,
(	847	)	,
(	846	)	,
(	846	)	,
(	845	)	,
(	845	)	,
(	844	)	,
(	844	)	,
(	843	)	,
(	842	)	,
(	842	)	,
(	841	)	,
(	841	)	,
(	840	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	838	)	,
(	837	)	,
(	836	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	834	)	,
(	833	)	,
(	833	)	,
(	832	)	,
(	832	)	,
(	831	)	,
(	830	)	,
(	830	)	,
(	829	)	,
(	829	)	,
(	828	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	823	)	,
(	823	)	,
(	822	)	,
(	822	)	,
(	821	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	819	)	,
(	818	)	,
(	817	)	,
(	817	)	,
(	816	)	,
(	816	)	,
(	815	)	,
(	815	)	,
(	814	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	811	)	,
(	811	)	,
(	810	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	808	)	,
(	807	)	,
(	807	)	,
(	806	)	,
(	805	)	,
(	805	)	,
(	804	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	797	)	,
(	796	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	793	)	,
(	793	)	,
(	792	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	785	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	775	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	755	)	,
(	754	)	,
(	754	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	748	)	,
(	748	)	,
(	747	)	,
(	747	)	,
(	746	)	,
(	746	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	741	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	736	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	730	)	,
(	730	)	,
(	729	)	,
(	729	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	700	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	697	)	,
(	696	)	,
(	695	)	,
(	695	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	692	)	,
(	691	)	,
(	690	)	,
(	690	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	683	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	666	)	,
(	666	)	,
(	665	)	,
(	664	)	,
(	664	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	661	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	655	)	,
(	655	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	650	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	646	)	,
(	646	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	642	)	,
(	642	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	626	)	,
(	626	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	622	)	,
(	622	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	616	)	,
(	616	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	610	)	,
(	610	)	,
(	609	)	,
(	608	)	,
(	608	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	598	)	,
(	598	)	,
(	597	)	,
(	596	)	,
(	595	)	,
(	595	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	591	)	,
(	591	)	,
(	590	)	,
(	589	)	,
(	589	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	574	)	,
(	574	)	,
(	573	)	,
(	572	)	,
(	572	)	,
(	571	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	567	)	,
(	567	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	561	)	,
(	561	)	,
(	560	)	,
(	559	)	,
(	558	)	,
(	558	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	523	)	,
(	523	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	508	)	,
(	508	)	,
(	507	)	,
(	506	)	,
(	505	)	,
(	505	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	482	)	,
(	482	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	478	)	,
(	478	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	461	)	,
(	461	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	457	)	,
(	457	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	447	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	443	)	,
(	443	)	,
(	442	)	,
(	441	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	432	)	,
(	431	)	,
(	430	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	427	)	,
(	427	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	415	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	409	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	399	)	,
(	398	)	,
(	397	)	,
(	397	)	,
(	396	)	,
(	396	)	,
(	395	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	393	)	,
(	393	)	,
(	392	)	,
(	392	)	,
(	391	)	,
(	391	)	,
(	390	)	,
(	390	)	,
(	389	)	,
(	388	)	,
(	388	)	,
(	387	)	,
(	387	)	,
(	386	)	,
(	386	)	,
(	385	)	,
(	385	)	,
(	384	)	,
(	384	)	,
(	383	)	,
(	383	)	,
(	382	)	,
(	382	)	,
(	381	)	,
(	381	)	,
(	380	)	,
(	380	)	,
(	380	)	,
(	379	)	,
(	379	)	,
(	378	)	,
(	378	)	,
(	377	)	,
(	377	)	,
(	376	)	,
(	376	)	,
(	375	)	,
(	375	)	,
(	374	)	,
(	374	)	,
(	373	)	,
(	373	)	,
(	372	)	,
(	372	)	,
(	372	)	,
(	371	)	,
(	371	)	,
(	370	)	,
(	370	)	,
(	369	)	,
(	369	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	367	)	,
(	367	)	,
(	366	)	,
(	366	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	364	)	,
(	364	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	362	)	,
(	362	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	360	)	,
(	360	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	358	)	,
(	358	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	355	)	,
(	355	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	347	)	,
(	347	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	349	)	,
(	349	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	351	)	,
(	351	)	,
(	352	)	,
(	352	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	354	)	,
(	354	)	,
(	355	)	,
(	355	)	,
(	356	)	,
(	356	)	,
(	357	)	,
(	357	)	,
(	358	)	,
(	358	)	,
(	359	)	,
(	359	)	,
(	360	)	,
(	360	)	,
(	361	)	,
(	361	)	,
(	362	)	,
(	362	)	,
(	363	)	,
(	364	)	,
(	364	)	,
(	365	)	,
(	365	)	,
(	366	)	,
(	366	)	,
(	367	)	,
(	368	)	,
(	368	)	,
(	369	)	,
(	369	)	,
(	370	)	,
(	371	)	,
(	371	)	,
(	372	)	,
(	373	)	,
(	373	)	,
(	374	)	,
(	375	)	,
(	375	)	,
(	376	)	,
(	377	)	,
(	377	)	,
(	378	)	,
(	379	)	,
(	379	)	,
(	380	)	,
(	381	)	,
(	381	)	,
(	382	)	,
(	383	)	,
(	384	)	,
(	384	)	,
(	385	)	,
(	386	)	,
(	387	)	,
(	387	)	,
(	388	)	,
(	389	)	,
(	390	)	,
(	390	)	,
(	391	)	,
(	392	)	,
(	393	)	,
(	394	)	,
(	394	)	,
(	395	)	,
(	396	)	,
(	397	)	,
(	398	)	,
(	399	)	,
(	399	)	,
(	400	)	,
(	401	)	,
(	402	)	,
(	403	)	,
(	404	)	,
(	405	)	,
(	406	)	,
(	406	)	,
(	407	)	,
(	408	)	,
(	409	)	,
(	410	)	,
(	411	)	,
(	412	)	,
(	413	)	,
(	414	)	,
(	415	)	,
(	416	)	,
(	417	)	,
(	418	)	,
(	419	)	,
(	420	)	,
(	421	)	,
(	422	)	,
(	423	)	,
(	424	)	,
(	425	)	,
(	426	)	,
(	427	)	,
(	428	)	,
(	429	)	,
(	430	)	,
(	431	)	,
(	432	)	,
(	433	)	,
(	434	)	,
(	435	)	,
(	437	)	,
(	438	)	,
(	439	)	,
(	440	)	,
(	441	)	,
(	442	)	,
(	443	)	,
(	444	)	,
(	446	)	,
(	447	)	,
(	448	)	,
(	449	)	,
(	450	)	,
(	451	)	,
(	453	)	,
(	454	)	,
(	455	)	,
(	456	)	,
(	457	)	,
(	459	)	,
(	460	)	,
(	461	)	,
(	462	)	,
(	464	)	,
(	465	)	,
(	466	)	,
(	467	)	,
(	469	)	,
(	470	)	,
(	471	)	,
(	473	)	,
(	474	)	,
(	475	)	,
(	477	)	,
(	478	)	,
(	479	)	,
(	481	)	,
(	482	)	,
(	483	)	,
(	485	)	,
(	486	)	,
(	488	)	,
(	489	)	,
(	490	)	,
(	492	)	,
(	493	)	,
(	495	)	,
(	496	)	,
(	497	)	,
(	499	)	,
(	500	)	,
(	502	)	,
(	503	)	,
(	505	)	,
(	506	)	,
(	508	)	,
(	509	)	,
(	511	)	,
(	512	)	,
(	514	)	,
(	515	)	,
(	517	)	,
(	518	)	,
(	520	)	,
(	522	)	,
(	523	)	,
(	525	)	,
(	526	)	,
(	528	)	,
(	530	)	,
(	531	)	,
(	533	)	,
(	534	)	,
(	536	)	,
(	538	)	,
(	539	)	,
(	541	)	,
(	543	)	,
(	544	)	,
(	546	)	,
(	548	)	,
(	549	)	,
(	551	)	,
(	553	)	,
(	555	)	,
(	556	)	,
(	558	)	,
(	560	)	,
(	562	)	,
(	563	)	,
(	565	)	,
(	567	)	,
(	569	)	,
(	570	)	,
(	572	)	,
(	574	)	,
(	576	)	,
(	578	)	,
(	580	)	,
(	581	)	,
(	583	)	,
(	585	)	,
(	587	)	,
(	589	)	,
(	591	)	,
(	593	)	,
(	595	)	,
(	597	)	,
(	598	)	,
(	600	)	,
(	602	)	,
(	604	)	,
(	606	)	,
(	608	)	,
(	610	)	,
(	612	)	,
(	614	)	,
(	616	)	,
(	618	)	,
(	620	)	,
(	622	)	,
(	624	)	,
(	626	)	,
(	628	)	,
(	630	)	,
(	633	)	,
(	635	)	,
(	637	)	,
(	639	)	,
(	641	)	,
(	643	)	,
(	645	)	,
(	647	)	,
(	650	)	,
(	652	)	,
(	654	)	,
(	656	)	,
(	658	)	,
(	660	)	,
(	663	)	,
(	665	)	,
(	667	)	,
(	669	)	,
(	672	)	,
(	674	)	,
(	676	)	,
(	678	)	,
(	681	)	,
(	683	)	,
(	685	)	,
(	687	)	,
(	690	)	,
(	692	)	,
(	694	)	,
(	697	)	,
(	699	)	,
(	701	)	,
(	704	)	,
(	706	)	,
(	709	)	,
(	711	)	,
(	713	)	,
(	716	)	,
(	718	)	,
(	721	)	,
(	723	)	,
(	726	)	,
(	728	)	,
(	731	)	,
(	733	)	,
(	736	)	,
(	738	)	,
(	741	)	,
(	743	)	,
(	746	)	,
(	748	)	,
(	751	)	,
(	753	)	,
(	756	)	,
(	759	)	,
(	761	)	,
(	764	)	,
(	766	)	,
(	769	)	,
(	772	)	,
(	774	)	,
(	777	)	,
(	780	)	,
(	782	)	,
(	785	)	,
(	788	)	,
(	790	)	,
(	793	)	,
(	796	)	,
(	799	)	,
(	801	)	,
(	804	)	,
(	807	)	,
(	810	)	,
(	812	)	,
(	815	)	,
(	818	)	,
(	821	)	,
(	824	)	,
(	827	)	,
(	829	)	,
(	832	)	,
(	835	)	,
(	838	)	,
(	841	)	,
(	844	)	,
(	847	)	,
(	850	)	,
(	853	)	,
(	856	)	,
(	859	)	,
(	861	)	,
(	864	)	,
(	867	)	,
(	870	)	,
(	873	)	,
(	877	)	,
(	880	)	,
(	883	)	,
(	886	)	,
(	889	)	,
(	892	)	,
(	895	)	,
(	898	)	,
(	901	)	,
(	904	)	,
(	907	)	,
(	911	)	,
(	914	)	,
(	917	)	,
(	920	)	,
(	923	)	,
(	926	)	,
(	930	)	,
(	933	)	,
(	936	)	,
(	939	)	,
(	943	)	,
(	946	)	,
(	949	)	,
(	952	)	,
(	956	)	,
(	959	)	,
(	962	)	,
(	966	)	,
(	969	)	,
(	972	)	,
(	976	)	,
(	979	)	,
(	983	)	,
(	986	)	,
(	989	)	,
(	993	)	,
(	996	)	,
(	1000	)	,
(	1003	)	,
(	1007	)	,
(	1010	)	,
(	1014	)	,
(	1017	)	,
(	1021	)	,
(	1024	)	,
(	1028	)	,
(	1031	)	,
(	1035	)	,
(	1038	)	,
(	1042	)	,
(	1046	)	,
(	1049	)	,
(	1053	)	,
(	1057	)	,
(	1060	)	,
(	1064	)	,
(	1068	)	,
(	1071	)	,
(	1075	)	,
(	1079	)	,
(	1082	)	,
(	1086	)	,
(	1090	)	,
(	1094	)	,
(	1097	)	,
(	1101	)	,
(	1105	)	,
(	1109	)	,
(	1113	)	,
(	1116	)	,
(	1120	)	,
(	1124	)	,
(	1128	)	,
(	1132	)	,
(	1136	)	,
(	1140	)	,
(	1144	)	,
(	1148	)	,
(	1152	)	,
(	1155	)	,
(	1159	)	,
(	1163	)	,
(	1167	)	,
(	1171	)	,
(	1175	)	,
(	1179	)	,
(	1184	)	,
(	1188	)	,
(	1192	)	,
(	1196	)	,
(	1200	)	,
(	1204	)	,
(	1208	)	,
(	1212	)	,
(	1216	)	,
(	1221	)	,
(	1225	)	,
(	1229	)	,
(	1233	)	,
(	1237	)	,
(	1242	)	,
(	1246	)	,
(	1250	)	,
(	1254	)	,
(	1259	)	,
(	1263	)	,
(	1267	)	,
(	1272	)	,
(	1276	)	,
(	1280	)	,
(	1285	)	,
(	1289	)	,
(	1293	)	,
(	1298	)	,
(	1302	)	,
(	1307	)	,
(	1311	)	,
(	1315	)	,
(	1320	)	,
(	1324	)	,
(	1329	)	,
(	1333	)	,
(	1338	)	,
(	1342	)	,
(	1347	)	,
(	1352	)	,
(	1356	)	,
(	1361	)	,
(	1365	)	,
(	1370	)	,
(	1375	)	,
(	1379	)	,
(	1384	)	,
(	1388	)	,
(	1393	)	,
(	1398	)	,
(	1403	)	,
(	1407	)	,
(	1412	)	,
(	1417	)	,
(	1422	)	,
(	1426	)	,
(	1431	)	,
(	1436	)	,
(	1441	)	,
(	1446	)	,
(	1450	)	,
(	1455	)	,
(	1460	)	,
(	1465	)	,
(	1470	)	,
(	1475	)	,
(	1480	)	,
(	1485	)	,
(	1490	)	,
(	1495	)	,
(	1500	)	,
(	1505	)	,
(	1510	)	,
(	1515	)	,
(	1520	)	,
(	1525	)	,
(	1530	)	,
(	1535	)	,
(	1540	)	,
(	1545	)	,
(	1550	)	,
(	1556	)	,
(	1561	)	,
(	1566	)	,
(	1571	)	,
(	1576	)	,
(	1581	)	,
(	1587	)	,
(	1592	)	,
(	1597	)	,
(	1603	)	,
(	1608	)	,
(	1613	)	,
(	1618	)	,
(	1624	)	,
(	1629	)	,
(	1635	)	,
(	1640	)	,
(	1645	)	,
(	1651	)	,
(	1656	)	,
(	1662	)	,
(	1667	)	,
(	1673	)	,
(	1678	)	,
(	1684	)	,
(	1689	)	,
(	1695	)	,
(	1700	)	,
(	1706	)	,
(	1711	)	,
(	1717	)	,
(	1722	)	,
(	1728	)	,
(	1734	)	,
(	1739	)	,
(	1745	)	,
(	1751	)	,
(	1756	)	,
(	1762	)	,
(	1768	)	,
(	1774	)	,
(	1779	)	,
(	1785	)	,
(	1791	)	,
(	1797	)	,
(	1803	)	,
(	1808	)	,
(	1814	)	,
(	1820	)	,
(	1826	)	,
(	1832	)	,
(	1838	)	,
(	1844	)	,
(	1850	)	,
(	1856	)	,
(	1862	)	,
(	1868	)	,
(	1874	)	,
(	1880	)	,
(	1886	)	,
(	1892	)	,
(	1898	)	,
(	1904	)	,
(	1910	)	,
(	1916	)	,
(	1922	)	,
(	1929	)	,
(	1935	)	,
(	1941	)	,
(	1947	)	,
(	1953	)	,
(	1960	)	,
(	1966	)	,
(	1972	)	,
(	1979	)	,
(	1985	)	,
(	1991	)	,
(	1997	)	,
(	2004	)	,
(	2010	)	,
(	2017	)	,
(	2023	)	,
(	2029	)	,
(	2036	)	,
(	2042	)	,
(	2049	)	,
(	2055	)	,
(	2062	)	,
(	2068	)	,
(	2075	)	,
(	2081	)	,
(	2088	)	,
(	2095	)	,
(	2101	)	,
(	2108	)	,
(	2114	)	,
(	2121	)	,
(	2128	)	,
(	2134	)	,
(	2141	)	,
(	2148	)	,
(	2155	)	,
(	2161	)	,
(	2168	)	,
(	2175	)	,
(	2182	)	,
(	2189	)	,
(	2195	)	,
(	2202	)	,
(	2209	)	,
(	2216	)	,
(	2223	)	,
(	2230	)	,
(	2237	)	,
(	2244	)	,
(	2251	)	,
(	2258	)	,
(	2265	)	,
(	2272	)	,
(	2279	)	,
(	2286	)	,
(	2293	)	,
(	2300	)	,
(	2307	)	,
(	2314	)	,
(	2321	)	,
(	2329	)	,
(	2336	)	,
(	2343	)	,
(	2350	)	,
(	2358	)	,
(	2365	)	,
(	2372	)	,
(	2379	)	,
(	2387	)	,
(	2394	)	,
(	2401	)	,
(	2409	)	,
(	2416	)	,
(	2424	)	,
(	2431	)	,
(	2438	)	,
(	2446	)	,
(	2453	)	,
(	2461	)	,
(	2468	)	,
(	2476	)	,
(	2483	)	,
(	2491	)	,
(	2499	)	,
(	2506	)	,
(	2514	)	,
(	2521	)	,
(	2529	)	,
(	2537	)	,
(	2544	)	,
(	2552	)	,
(	2560	)	,
(	2568	)	,
(	2575	)	,
(	2583	)	,
(	2591	)	,
(	2599	)	,
(	2607	)	,
(	2615	)	,
(	2622	)	,
(	2630	)	,
(	2638	)	,
(	2646	)	,
(	2654	)	,
(	2662	)	,
(	2670	)	,
(	2678	)	,
(	2686	)	,
(	2694	)	,
(	2702	)	,
(	2710	)	,
(	2718	)	,
(	2727	)	,
(	2735	)	,
(	2743	)	,
(	2751	)	,
(	2759	)	,
(	2767	)	,
(	2776	)	,
(	2784	)	,
(	2792	)	,
(	2801	)	,
(	2809	)	,
(	2817	)	,
(	2826	)	,
(	2834	)	,
(	2842	)	,
(	2851	)	,
(	2859	)	,
(	2868	)	,
(	2876	)	,
(	2885	)	,
(	2893	)	,
(	2902	)	,
(	2910	)	,
(	2919	)	,
(	2927	)	,
(	2936	)	,
(	2945	)	,
(	2953	)	,
(	2962	)	,
(	2971	)	,
(	2979	)	,
(	2988	)	,
(	2997	)	,
(	3006	)	,
(	3014	)	,
(	3023	)	,
(	3032	)	,
(	3041	)	,
(	3050	)	,
(	3059	)	,
(	3067	)	,
(	3076	)	,
(	3085	)	,
(	3094	)	,
(	3103	)	,
(	3112	)	,
(	3121	)	,
(	3130	)	,
(	3139	)	,
(	3149	)	,
(	3158	)	,
(	3167	)	,
(	3176	)	,
(	3185	)	,
(	3194	)	,
(	3203	)	,
(	3213	)	,
(	3222	)	,
(	3231	)	,
(	3241	)	,
(	3250	)	,
(	3259	)	,
(	3269	)	,
(	3278	)	,
(	3287	)	,
(	3297	)	,
(	3306	)	,
(	3316	)	,
(	3325	)	,
(	3335	)	,
(	3344	)	,
(	3354	)	,
(	3363	)	,
(	3373	)	,
(	3382	)	,
(	3392	)	,
(	3402	)	,
(	3411	)	,
(	3421	)	,
(	3431	)	,
(	3441	)	,
(	3450	)	,
(	3460	)	,
(	3470	)	,
(	3480	)	,
(	3490	)	,
(	3499	)	,
(	3509	)	,
(	3519	)	,
(	3529	)	,
(	3539	)	,
(	3549	)	,
(	3559	)	,
(	3569	)	,
(	3579	)	,
(	3589	)	,
(	3599	)	,
(	3609	)	,
(	3619	)	,
(	3630	)	,
(	3640	)	,
(	3650	)	,
(	3660	)	,
(	3670	)	,
(	3681	)	,
(	3691	)	,
(	3701	)	,
(	3711	)	,
(	3722	)	,
(	3732	)	,
(	3743	)	,
(	3753	)	,
(	3763	)	,
(	3774	)	,
(	3784	)	,
(	3795	)	,
(	3805	)	,
(	3816	)	,
(	3826	)	,
(	3837	)	,
(	3848	)	,
(	3858	)	,
(	3869	)	,
(	3880	)	,
(	3890	)	,
(	3901	)	,
(	3912	)	,
(	3922	)	,
(	3933	)	,
(	3944	)	,
(	3955	)	,
(	3966	)	,
(	3977	)	,
(	3988	)	,
(	3998	)	,
(	4009	)	,
(	4020	)	,
(	4031	)	,
(	4042	)	,
(	4053	)	,
(	4064	)	,
(	4076	)	,
(	4087	)	,
(	4098	)	,
(	4109	)	,
(	4120	)	,
(	4131	)	,
(	4142	)	,
(	4154	)	,
(	4165	)	,
(	4176	)	,
(	4188	)	,
(	4199	)	,
(	4210	)	,
(	4222	)	,
(	4233	)	,
(	4245	)	,
(	4256	)	,
(	4267	)	,
(	4279	)	,
(	4290	)	,
(	4302	)	,
(	4314	)	,
(	4325	)	,
(	4337	)	,
(	4348	)	,
(	4360	)	,
(	4372	)	,
(	4383	)	,
(	4395	)	,
(	4407	)	,
(	4419	)	,
(	4431	)	,
(	4442	)	,
(	4454	)	,
(	4466	)	,
(	4478	)	,
(	4490	)	,
(	4502	)	,
(	4514	)	,
(	4526	)	,
(	4538	)	,
(	4550	)	,
(	4562	)	,
(	4574	)	,
(	4586	)	,
(	4598	)	,
(	4611	)	,
(	4623	)	,
(	4635	)	,
(	4647	)	,
(	4659	)	,
(	4672	)	,
(	4684	)	,
(	4696	)	,
(	4709	)	,
(	4721	)	,
(	4734	)	,
(	4746	)	,
(	4759	)	,
(	4771	)	,
(	4784	)	,
(	4796	)	,
(	4809	)	,
(	4821	)	,
(	4834	)	,
(	4846	)	,
(	4859	)	,
(	4872	)	,
(	4885	)	,
(	4897	)	,
(	4910	)	,
(	4923	)	,
(	4936	)	,
(	4948	)	,
(	4961	)	,
(	4974	)	,
(	4987	)	,
(	5000	)	,
(	5013	)	,
(	5026	)	,
(	5039	)	,
(	5052	)	,
(	5065	)	,
(	5078	)	,
(	5091	)	,
(	5104	)	,
(	5118	)	,
(	5131	)	,
(	5144	)	,
(	5157	)	,
(	5171	)	,
(	5184	)	,
(	5197	)	,
(	5211	)	,
(	5224	)	,
(	5237	)	,
(	5251	)	,
(	5264	)	,
(	5278	)	,
(	5291	)	,
(	5305	)	,
(	5318	)	,
(	5332	)	,
(	5345	)	,
(	5359	)	,
(	5373	)	,
(	5386	)	,
(	5400	)	,
(	5414	)	,
(	5428	)	,
(	5441	)	,
(	5455	)	,
(	5469	)	,
(	5483	)	,
(	5497	)	,
(	5511	)	,
(	5525	)	,
(	5539	)	,
(	5553	)	,
(	5567	)	,
(	5581	)	,
(	5595	)	,
(	5609	)	,
(	5623	)	,
(	5637	)	,
(	5651	)	,
(	5666	)	,
(	5680	)	,
(	5694	)	,
(	5709	)	,
(	5723	)	,
(	5737	)	,
(	5752	)	,
(	5766	)	,
(	5780	)	,
(	5795	)	,
(	5809	)	,
(	5824	)	,
(	5838	)	,
(	5853	)	,
(	5868	)	,
(	5882	)	,
(	5897	)	,
(	5912	)	,
(	5926	)	,
(	5941	)	,
(	5956	)	,
(	5970	)	,
(	5985	)	,
(	6000	)	,
(	6015	)	,
(	6030	)	,
(	6045	)	,
(	6060	)	,
(	6075	)	,
(	6090	)	,
(	6105	)	,
(	6120	)	,
(	6135	)	,
(	6150	)	,
(	6165	)	,
(	6180	)	,
(	6196	)	,
(	6211	)	,
(	6226	)	,
(	6241	)	,
(	6257	)	,
(	6272	)	,
(	6287	)	,
(	6303	)	,
(	6318	)	,
(	6334	)	,
(	6349	)	,
(	6365	)	,
(	6380	)	,
(	6396	)	,
(	6411	)	,
(	6427	)	,
(	6443	)	,
(	6458	)	,
(	6474	)	,
(	6490	)	,
(	6506	)	,
(	6521	)	,
(	6537	)	,
(	6553	)	,
(	6569	)	,
(	6585	)	,
(	6601	)	,
(	6617	)	,
(	6633	)	,
(	6649	)	,
(	6665	)	,
(	6681	)	,
(	6697	)	,
(	6713	)	,
(	6729	)	,
(	6746	)	,
(	6762	)	,
(	6778	)	,
(	6794	)	,
(	6811	)	,
(	6827	)	,
(	6843	)	,
(	6860	)	,
(	6876	)	,
(	6893	)	,
(	6909	)	,
(	6926	)	,
(	6942	)	,
(	6959	)	,
(	6975	)	,
(	6992	)	,
(	7009	)	,
(	7025	)	,
(	7042	)	,
(	7059	)	,
(	7076	)	,
(	7093	)	,
(	7109	)	,
(	7126	)	,
(	7143	)	,
(	7160	)	,
(	7177	)	,
(	7194	)	,
(	7211	)	,
(	7228	)	,
(	7245	)	,
(	7262	)	,
(	7280	)	,
(	7297	)	,
(	7314	)	,
(	7331	)	,
(	7349	)	,
(	7366	)	,
(	7383	)	,
(	7401	)	,
(	7418	)	,
(	7435	)	,
(	7453	)	,
(	7470	)	,
(	7488	)	,
(	7505	)	,
(	7523	)	,
(	7541	)	,
(	7558	)	,
(	7576	)	,
(	7594	)	,
(	7611	)	,
(	7629	)	,
(	7647	)	,
(	7665	)	,
(	7683	)	,
(	7700	)	,
(	7718	)	,
(	7736	)	,
(	7754	)	,
(	7772	)	,
(	7790	)	,
(	7808	)	,
(	7826	)	,
(	7845	)	,
(	7863	)	,
(	7881	)	,
(	7899	)	,
(	7917	)	,
(	7936	)	,
(	7954	)	,
(	7972	)	,
(	7991	)	,
(	8009	)	,
(	8028	)	,
(	8046	)	,
(	8065	)	,
(	8083	)	,
(	8102	)	,
(	8120	)	,
(	8139	)	,
(	8158	)	,
(	8176	)	,
(	8195	)	,
(	8214	)	,
(	8233	)	,
(	8252	)	,
(	8270	)	,
(	8289	)	,
(	8308	)	,
(	8327	)	,
(	8346	)	,
(	8365	)	,
(	8384	)	,
(	8403	)	,
(	8423	)	,
(	8442	)	,
(	8461	)	,
(	8480	)	,
(	8499	)	,
(	8519	)	,
(	8538	)	,
(	8557	)	,
(	8577	)	,
(	8596	)	,
(	8616	)	,
(	8635	)	,
(	8655	)	,
(	8674	)	,
(	8694	)	,
(	8713	)	,
(	8733	)	,
(	8753	)	,
(	8772	)	,
(	8792	)	,
(	8812	)	,
(	8832	)	,
(	8851	)	,
(	8871	)	,
(	8891	)	,
(	8911	)	,
(	8931	)	,
(	8951	)	,
(	8971	)	,
(	8991	)	,
(	9011	)	,
(	9032	)	,
(	9052	)	,
(	9072	)	,
(	9092	)	,
(	9112	)	,
(	9133	)	,
(	9153	)	,
(	9173	)	,
(	9194	)	,
(	9214	)	,
(	9235	)	,
(	9255	)	,
(	9276	)	,
(	9296	)	,
(	9317	)	,
(	9338	)	,
(	9358	)	,
(	9379	)	,
(	9400	)	,
(	9421	)	,
(	9441	)	,
(	9462	)	,
(	9483	)	,
(	9504	)	,
(	9525	)	,
(	9546	)	,
(	9567	)	,
(	9588	)	,
(	9609	)	,
(	9630	)	,
(	9651	)	,
(	9673	)	,
(	9694	)	,
(	9715	)	,
(	9736	)	,
(	9758	)	,
(	9779	)	,
(	9801	)	,
(	9822	)	,
(	9843	)	,
(	9865	)	,
(	9887	)	,
(	9908	)	,
(	9930	)	,
(	9951	)	,
(	9973	)	,
(	9995	)	,
(	10017	)	,
(	10038	)	,
(	10060	)	,
(	10082	)	,
(	10104	)	,
(	10126	)	,
(	10148	)	,
(	10170	)	,
(	10192	)	,
(	10214	)	,
(	10236	)	,
(	10258	)	,
(	10280	)	,
(	10303	)	,
(	10325	)	,
(	10347	)	,
(	10369	)	,
(	10392	)	,
(	10414	)	,
(	10437	)	,
(	10459	)	,
(	10482	)	,
(	10504	)	,
(	10527	)	,
(	10549	)	,
(	10572	)	,
(	10595	)	,
(	10617	)	,
(	10640	)	,
(	10663	)	,
(	10686	)	,
(	10709	)	,
(	10731	)	,
(	10754	)	,
(	10777	)	,
(	10800	)	,
(	10823	)	,
(	10846	)	,
(	10870	)	,
(	10893	)	,
(	10916	)	,
(	10939	)	,
(	10962	)	,
(	10986	)	,
(	11009	)	,
(	11032	)	,
(	11056	)	,
(	11079	)	,
(	11103	)	,
(	11126	)	,
(	11150	)	,
(	11173	)	,
(	11197	)	,
(	11221	)	,
(	11244	)	,
(	11268	)	,
(	11292	)	,
(	11316	)	,
(	11340	)	,
(	11363	)	,
(	11387	)	,
(	11411	)	,
(	11435	)	,
(	11459	)	,
(	11483	)	,
(	11508	)	,
(	11532	)	,
(	11556	)	,
(	11580	)	,
(	11604	)	,
(	11629	)	,
(	11653	)	,
(	11677	)	,
(	11702	)	,
(	11726	)	,
(	11751	)	,
(	11775	)	,
(	11800	)	,
(	11824	)	,
(	11849	)	,
(	11874	)	,
(	11899	)	,
(	11923	)	,
(	11948	)	,
(	11973	)	,
(	11998	)	,
(	12023	)	,
(	12048	)	,
(	12073	)	,
(	12098	)	,
(	12123	)	,
(	12148	)	,
(	12173	)	,
(	12198	)	,
(	12223	)	,
(	12249	)	,
(	12274	)	,
(	12299	)	,
(	12325	)	,
(	12350	)	,
(	12375	)	,
(	12401	)	,
(	12426	)	,
(	12452	)	,
(	12478	)	,
(	12503	)	,
(	12529	)	,
(	12555	)	,
(	12580	)	,
(	12606	)	,
(	12632	)	,
(	12658	)	,
(	12684	)	,
(	12710	)	,
(	12736	)	,
(	12762	)	,
(	12788	)	,
(	12814	)	,
(	12840	)	,
(	12866	)	,
(	12893	)	,
(	12919	)	,
(	12945	)	,
(	12972	)	,
(	12998	)	,
(	13024	)	,
(	13051	)	,
(	13077	)	,
(	13104	)	,
(	13131	)	,
(	13157	)	,
(	13184	)	,
(	13211	)	,
(	13237	)	,
(	13264	)	,
(	13291	)	,
(	13318	)	,
(	13345	)	,
(	13372	)	,
(	13399	)	,
(	13426	)	,
(	13453	)	,
(	13480	)	,
(	13507	)	,
(	13534	)	,
(	13562	)	,
(	13589	)	,
(	13616	)	,
(	13644	)	,
(	13671	)	,
(	13698	)	,
(	13726	)	,
(	13753	)	,
(	13781	)	,
(	13809	)	,
(	13836	)	,
(	13864	)	,
(	13892	)	,
(	13919	)	,
(	13947	)	,
(	13975	)	,
(	14003	)	,
(	14031	)	,
(	14059	)	,
(	14087	)	,
(	14115	)	,
(	14143	)	,
(	14171	)	,
(	14199	)	,
(	14228	)	,
(	14256	)	,
(	14284	)	,
(	14312	)	,
(	14341	)	,
(	14369	)	,
(	14398	)	,
(	14426	)	,
(	14455	)	,
(	14483	)	,
(	14512	)	,
(	14541	)	,
(	14569	)	,
(	14598	)	,
(	14627	)	,
(	14656	)	,
(	14685	)	,
(	14714	)	,
(	14743	)	,
(	14772	)	,
(	14801	)	,
(	14830	)	,
(	14859	)	,
(	14888	)	,
(	14917	)	,
(	14947	)	,
(	14976	)	,
(	15005	)	,
(	15035	)	,
(	15064	)	,
(	15094	)	,
(	15123	)	,
(	15153	)	,
(	15182	)	,
(	15212	)	,
(	15242	)	,
(	15272	)	,
(	15301	)	,
(	15331	)	,
(	15361	)	,
(	15391	)	,
(	15421	)	,
(	15451	)	,
(	15481	)	,
(	15511	)	,
(	15541	)	,
(	15571	)	,
(	15602	)	,
(	15632	)	,
(	15662	)	,
(	15692	)	,
(	15723	)	,
(	15753	)	,
(	15784	)	,
(	15814	)	,
(	15845	)	,
(	15875	)	,
(	15906	)	,
(	15937	)	,
(	15968	)	,
(	15998	)	,
(	16029	)	,
(	16060	)	,
(	16091	)	,
(	16122	)	,
(	16153	)	,
(	16184	)	,
(	16215	)	,
(	16246	)	,
(	16277	)	,
(	16309	)	,
(	16340	)	,
(	16371	)	,
(	16403	)	,
(	16434	)	,
(	16465	)	,
(	16497	)	,
(	16528	)	,
(	16560	)	,
(	16592	)	,
(	16623	)	,
(	16655	)	,
(	16687	)	,
(	16719	)	,
(	16750	)	,
(	16782	)	,
(	16814	)	,
(	16846	)	,
(	16878	)	,
(	16910	)	,
(	16943	)	,
(	16975	)	,
(	17007	)	,
(	17039	)	,
(	17071	)	,
(	17104	)	,
(	17136	)	,
(	17169	)	,
(	17201	)	,
(	17234	)	,
(	17266	)	,
(	17299	)	,
(	17332	)	,
(	17364	)	,
(	17397	)	,
(	17430	)	,
(	17463	)	,
(	17496	)	,
(	17528	)	,
(	17561	)	,
(	17595	)	,
(	17628	)	,
(	17661	)	,
(	17694	)	,
(	17727	)	,
(	17760	)	,
(	17794	)	,
(	17827	)	,
(	17860	)	,
(	17894	)	,
(	17927	)	,
(	17961	)	,
(	17994	)	,
(	18028	)	,
(	18062	)	,
(	18096	)	,
(	18129	)	,
(	18163	)	,
(	18197	)	,
(	18231	)	,
(	18265	)	,
(	18299	)	,
(	18333	)	,
(	18367	)	,
(	18401	)	,
(	18435	)	,
(	18470	)	,
(	18504	)	,
(	18538	)	,
(	18573	)	,
(	18607	)	,
(	18642	)	,
(	18676	)	,
(	18711	)	,
(	18745	)	,
(	18780	)	,
(	18815	)	,
(	18849	)	,
(	18884	)	,
(	18919	)	,
(	18954	)	,
(	18989	)	,
(	19024	)	,
(	19059	)	,
(	19094	)	,
(	19129	)	,
(	19164	)	,
(	19200	)	,
(	19235	)	,
(	19270	)	,
(	19306	)	,
(	19341	)	,
(	19377	)	,
(	19412	)	,
(	19448	)	,
(	19483	)	,
(	19519	)	,
(	19555	)	,
(	19590	)	,
(	19626	)	,
(	19662	)	,
(	19698	)	,
(	19734	)	,
(	19770	)	,
(	19806	)	,
(	19842	)	,
(	19878	)	,
(	19915	)	,
(	19951	)	,
(	19987	)	,
(	20023	)	,
(	20060	)	,
(	20096	)	,
(	20133	)	,
(	20169	)	,
(	20206	)	,
(	20243	)	,
(	20279	)	,
(	20316	)	,
(	20353	)	,
(	20390	)	,
(	20427	)	,
(	20464	)	,
(	20501	)	,
(	20538	)	,
(	20575	)	,
(	20612	)	,
(	20649	)	,
(	20686	)	,
(	20723	)	,
(	20761	)	,
(	20798	)	,
(	20836	)	,
(	20873	)	,
(	20911	)	,
(	20948	)	,
(	20986	)	,
(	21024	)	,
(	21061	)	,
(	21099	)	,
(	21137	)	,
(	21175	)	,
(	21213	)	,
(	21251	)	,
(	21289	)	,
(	21327	)	,
(	21365	)	,
(	21403	)	,
(	21442	)	,
(	21480	)	,
(	21518	)	,
(	21557	)	,
(	21595	)	,
(	21633	)	,
(	21672	)	,
(	21711	)	,
(	21749	)	,
(	21788	)	,
(	21827	)	,
(	21866	)	,
(	21904	)	,
(	21943	)	,
(	21982	)	,
(	22021	)	,
(	22060	)	,
(	22099	)	,
(	22139	)	,
(	22178	)	,
(	22217	)	,
(	22256	)	,
(	22296	)	,
(	22335	)	,
(	22375	)	,
(	22414	)	,
(	22454	)	,
(	22493	)	,
(	22533	)	,
(	22573	)	,
(	22612	)	,
(	22652	)	,
(	22692	)	,
(	22732	)	,
(	22772	)	,
(	22812	)	,
(	22852	)	,
(	22892	)	,
(	22933	)	,
(	22973	)	,
(	23013	)	,
(	23053	)	,
(	23094	)	,
(	23134	)	,
(	23175	)	,
(	23215	)	,
(	23256	)	,
(	23297	)	,
(	23337	)	,
(	23378	)	,
(	23419	)	,
(	23460	)	,
(	23501	)	,
(	23542	)	,
(	23583	)	,
(	23624	)	,
(	23665	)	,
(	23706	)	,
(	23747	)	,
(	23789	)	,
(	23830	)	,
(	23872	)	,
(	23913	)	,
(	23955	)	,
(	23996	)	,
(	24038	)	,
(	24079	)	,
(	24121	)	,
(	24163	)	,
(	24205	)	,
(	24247	)	,
(	24289	)	,
(	24331	)	,
(	24373	)	,
(	24415	)	,
(	24457	)	,
(	24499	)	,
(	24541	)	,
(	24584	)	,
(	24626	)	,
(	24668	)	,
(	24711	)	,
(	24753	)	,
(	24796	)	,
(	24839	)	,
(	24881	)	,
(	24924	)	,
(	24967	)	,
(	25010	)	,
(	25053	)	,
(	25096	)	,
(	25139	)	,
(	25182	)	,
(	25225	)	,
(	25268	)

);

end package LUT_pkg;
